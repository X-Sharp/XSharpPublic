#define abc "���"

