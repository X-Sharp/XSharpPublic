// test include file
#define XSharp TheBest