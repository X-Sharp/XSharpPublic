///////////////////////////////////////////////////////////////////////////
// VOSystemLibrary.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// System Classes library
//

#define SE_ABORT 0
#define SE_IGNORE 1
#define SE_RETRY 2
#define SE_CANCEL 3
#define SE_OK 4
#define SE_YES 5
#define SE_NO 6
#define SE_CLOSE 7
#define SE_DEFAULT 0x80000000
#define E_DEFAULT FALSE
#define E_RETRY TRUE
#define E_EXCEPTION 5333L
#define E_ACCESSVIOLATION (5333L)
#define E_DATATYPE_MISALIGNMENT (5334L)
#define E_SINGLE_STEP (5335L)
#define E_ARRAY_BOUNDS_EXCEEDED (5336L)
#define E_FLT_DENORMAL_OPERAND (5337L)
#define E_FLT_DIVIDE_BY_ZERO (5338L)
#define E_FLT_INEXACT_RESULT (5339L)
#define E_FLT_INVALID_OPERATION (5340L)
#define E_FLT_OVERFLOW (5341L)
#define E_FLT_STACK_CHECK (5342L)
#define E_FLT_UNDERFLOW (5343L)
#define E_INT_DIVIDE_BY_ZERO (5344L)
#define E_INT_OVERFLOW (5345L)
#define E_PRIV_INSTRUCTION (5346L)
#define E_ILLEGAL_INSTRUCTION (5347L)
#define E_NONCONTINUABLE_EXCEPTION (5348L)
#define E_STACK_OVERFLOW (5349L)
#define E_INVALID_DISPOSITION (5350L)
#define E_GUARD_PAGE (5351L)
#define EC_ALERT 0
#define EC_IGNORE 1
#define EC_RETRY 2
#define EC_BREAK 3
#define EG_APPENDLOCK 40
#define EG_ARG 1
#define EG_BADALIAS 17
#define EG_BADPAGEFAULT 52
#define EG_BADPTR 51
#define EG_BOUND 2
#define EG_CLOSE 22
#define EG_COMPLEXITY 8
#define EG_CORRUPTION 32
#define EG_CREATE 20
#define EG_DATATYPE 33
#define EG_DATAWIDTH 34
#define EG_DUPALIAS 18
#define EG_DYNPTR 54
#define EG_ERRORBLOCK 49
#define EG_ERRORBUILD 53
#define EG_EVALSTACK 48
#define EG_LIMIT 31
#define EG_LOCK 41
#define EG_LOCK_ERROR 45
#define EG_LOCK_TIMEOUT 46
#define EG_MEM 11
#define EG_MEMOVERFLOW 9
#define EG_NOALIAS 15
#define EG_NOATOM 26
#define EG_NOCLASS 27
#define EG_NOFUNC 12
#define EG_NOMETHOD 13
#define EG_NOORDER 36
#define EG_NOTABLE 35
#define EG_NOVAR 14
#define EG_NOVARMETHOD 16
#define EG_NUMERR 6
#define EG_NUMOVERFLOW 4
#define EG_OPEN 21
#define EG_PRINT 25
#define EG_PROTECTION 50
#define EG_READ 23
#define EG_READONLY 39
#define EG_REFERENCE 29
#define EG_SEQUENCE 10
#define EG_SHARED 37
#define EG_STACK 47
#define EG_STROVERFLOW 3
#define EG_SYNTAX 7
#define EG_UNLOCKED 38
#define EG_UNSUPPORTED 30
#define EG_WRITE 24
#define EG_WRONGCLASS 28
#define EG_ZERODIV 5
#define ES_CATASTROPHIC 3
#define ES_ERROR 2
#define ES_WARNING 1
#define ES_WHOCARES 0
#define REG_BUFF_SIZE 64
#define INT_WINDOWS 1
#define INT_CLIPPER 0
#define INT_BINARY 2
#define RT_MSG_MONTH 4095
#define RT_MSG_DAY 4107
#define RT_MSG_LITERAL 8192
#define RT_MSG_LITERAL_MAX 10
#define RT_MSG_DOSERR 16448
#define RT_MSG_MONTH1 (RT_MSG_MONTH + 1)
#define RT_MSG_MONTH2 (RT_MSG_MONTH + 2)
#define RT_MSG_MONTH3 (RT_MSG_MONTH + 3)
#define RT_MSG_MONTH4 (RT_MSG_MONTH + 4)
#define RT_MSG_MONTH5 (RT_MSG_MONTH + 5)
#define RT_MSG_MONTH6 (RT_MSG_MONTH + 6)
#define RT_MSG_MONTH7 (RT_MSG_MONTH + 7)
#define RT_MSG_MONTH8 (RT_MSG_MONTH + 8)
#define RT_MSG_MONTH9 (RT_MSG_MONTH + 9)
#define RT_MSG_MONTH10 (RT_MSG_MONTH + 10)
#define RT_MSG_MONTH11 (RT_MSG_MONTH + 11)
#define RT_MSG_MONTH12 (RT_MSG_MONTH + 12)
#define RT_MSG_DAY1 (RT_MSG_DAY + 1)
#define RT_MSG_DAY2 (RT_MSG_DAY + 2)
#define RT_MSG_DAY3 (RT_MSG_DAY + 3)
#define RT_MSG_DAY4 (RT_MSG_DAY + 4)
#define RT_MSG_DAY5 (RT_MSG_DAY + 5)
#define RT_MSG_DAY6 (RT_MSG_DAY + 6)
#define RT_MSG_DAY7 (RT_MSG_DAY + 7)
#define RT_MSG_INFOSTRING (4115)
#define RT_MSG_SHORT_TRUE (RT_MSG_LITERAL + 1)
#define RT_MSG_SHORT_FALSE (RT_MSG_LITERAL + 2)
#define RT_MSG_LONG_TRUE (RT_MSG_LITERAL + 3)
#define RT_MSG_LONG_FALSE (RT_MSG_LITERAL + 4)
#define RT_MSG_SHORT_YES (RT_MSG_LITERAL + 5)
#define RT_MSG_SHORT_NO (RT_MSG_LITERAL + 6)
#define RT_MSG_LONG_YES (RT_MSG_LITERAL + 7)
#define RT_MSG_LONG_NO (RT_MSG_LITERAL + 8)
#define RT_MSG_CURRENCY (RT_MSG_LITERAL + 9)
#define RT_MSG_YNSTRING (RT_MSG_LITERAL + 10)
#define RT_MSG_DOSERR_0 (RT_MSG_DOSERR + 0)
#define RT_MSG_DOSERR_1 (RT_MSG_DOSERR + 1)
#define RT_MSG_DOSERR_2 (RT_MSG_DOSERR + 2)
#define RT_MSG_DOSERR_3 (RT_MSG_DOSERR + 3)
#define RT_MSG_DOSERR_4 (RT_MSG_DOSERR + 4)
#define RT_MSG_DOSERR_5 (RT_MSG_DOSERR + 5)
#define RT_MSG_DOSERR_6 (RT_MSG_DOSERR + 6)
#define RT_MSG_DOSERR_7 (RT_MSG_DOSERR + 7)
#define RT_MSG_DOSERR_8 (RT_MSG_DOSERR + 8)
#define RT_MSG_DOSERR_9 (RT_MSG_DOSERR + 9)
#define RT_MSG_DOSERR_10 (RT_MSG_DOSERR + 10)
#define RT_MSG_DOSERR_11 (RT_MSG_DOSERR + 11)
#define RT_MSG_DOSERR_12 (RT_MSG_DOSERR + 12)
#define RT_MSG_DOSERR_13 (RT_MSG_DOSERR + 13)
#define RT_MSG_DOSERR_14 (RT_MSG_DOSERR + 14)
#define RT_MSG_DOSERR_15 (RT_MSG_DOSERR + 15)
#define RT_MSG_DOSERR_16 (RT_MSG_DOSERR + 16)
#define RT_MSG_DOSERR_17 (RT_MSG_DOSERR + 17)
#define RT_MSG_DOSERR_18 (RT_MSG_DOSERR + 18)
#define RT_MSG_DOSERR_19 (RT_MSG_DOSERR + 19)
#define RT_MSG_DOSERR_20 (RT_MSG_DOSERR + 20)
#define RT_MSG_DOSERR_21 (RT_MSG_DOSERR + 21)
#define RT_MSG_DOSERR_22 (RT_MSG_DOSERR + 22)
#define RT_MSG_DOSERR_23 (RT_MSG_DOSERR + 23)
#define RT_MSG_DOSERR_24 (RT_MSG_DOSERR + 24)
#define RT_MSG_DOSERR_25 (RT_MSG_DOSERR + 25)
#define RT_MSG_DOSERR_26 (RT_MSG_DOSERR + 26)
#define RT_MSG_DOSERR_27 (RT_MSG_DOSERR + 27)
#define RT_MSG_DOSERR_28 (RT_MSG_DOSERR + 28)
#define RT_MSG_DOSERR_29 (RT_MSG_DOSERR + 29)
#define RT_MSG_DOSERR_30 (RT_MSG_DOSERR + 30)
#define RT_MSG_DOSERR_31 (RT_MSG_DOSERR + 31)
#define RT_MSG_DOSERR_32 (RT_MSG_DOSERR + 32)
#define RT_MSG_DOSERR_33 (RT_MSG_DOSERR + 33)
#define RT_MSG_DOSERR_34 (RT_MSG_DOSERR + 34)
#define RT_MSG_DOSERR_35 (RT_MSG_DOSERR + 35)
#define RT_MSG_DOSERR_36 (RT_MSG_DOSERR + 36)
#define RT_MSG_DOSERR_37 (RT_MSG_DOSERR + 37)
#define RT_MSG_DOSERR_38 (RT_MSG_DOSERR + 38)
#define RT_MSG_DOSERR_39 (RT_MSG_DOSERR + 39)
#define RT_MSG_DOSERR_40 (RT_MSG_DOSERR + 40)
#define RT_MSG_DOSERR_41 (RT_MSG_DOSERR + 41)
#define RT_MSG_DOSERR_42 (RT_MSG_DOSERR + 42)
#define RT_MSG_DOSERR_43 (RT_MSG_DOSERR + 43)
#define RT_MSG_DOSERR_44 (RT_MSG_DOSERR + 44)
#define RT_MSG_DOSERR_45 (RT_MSG_DOSERR + 45)
#define RT_MSG_DOSERR_46 (RT_MSG_DOSERR + 46)
#define RT_MSG_DOSERR_47 (RT_MSG_DOSERR + 47)
#define RT_MSG_DOSERR_48 (RT_MSG_DOSERR + 48)
#define RT_MSG_DOSERR_49 (RT_MSG_DOSERR + 49)
#define RT_MSG_DOSERR_50 (RT_MSG_DOSERR + 50)
#define RT_MSG_DOSERR_51 (RT_MSG_DOSERR + 51)
#define RT_MSG_DOSERR_52 (RT_MSG_DOSERR + 52)
#define RT_MSG_DOSERR_53 (RT_MSG_DOSERR + 53)
#define RT_MSG_DOSERR_54 (RT_MSG_DOSERR + 54)
#define RT_MSG_DOSERR_55 (RT_MSG_DOSERR + 55)
#define RT_MSG_DOSERR_56 (RT_MSG_DOSERR + 56)
#define RT_MSG_DOSERR_57 (RT_MSG_DOSERR + 57)
#define RT_MSG_DOSERR_58 (RT_MSG_DOSERR + 58)
#define RT_MSG_DOSERR_59 (RT_MSG_DOSERR + 59)
#define RT_MSG_DOSERR_60 (RT_MSG_DOSERR + 60)
#define RT_MSG_DOSERR_61 (RT_MSG_DOSERR + 61)
#define RT_MSG_DOSERR_62 (RT_MSG_DOSERR + 62)
#define RT_MSG_DOSERR_63 (RT_MSG_DOSERR + 63)
#define RT_MSG_DOSERR_64 (RT_MSG_DOSERR + 64)
#define RT_MSG_DOSERR_65 (RT_MSG_DOSERR + 65)
#define RT_MSG_DOSERR_66 (RT_MSG_DOSERR + 66)
#define RT_MSG_DOSERR_67 (RT_MSG_DOSERR + 67)
#define RT_MSG_DOSERR_68 (RT_MSG_DOSERR + 68)
#define RT_MSG_DOSERR_69 (RT_MSG_DOSERR + 69)
#define RT_MSG_DOSERR_70 (RT_MSG_DOSERR + 70)
#define RT_MSG_DOSERR_71 (RT_MSG_DOSERR + 71)
#define RT_MSG_DOSERR_72 (RT_MSG_DOSERR + 72)
#define RT_MSG_DOSERR_73 (RT_MSG_DOSERR + 73)
#define RT_MSG_DOSERR_74 (RT_MSG_DOSERR + 74)
#define RT_MSG_DOSERR_75 (RT_MSG_DOSERR + 75)
#define RT_MSG_DOSERR_76 (RT_MSG_DOSERR + 76)
#define RT_MSG_DOSERR_77 (RT_MSG_DOSERR + 77)
#define RT_MSG_DOSERR_78 (RT_MSG_DOSERR + 78)
#define RT_MSG_DOSERR_79 (RT_MSG_DOSERR + 79)
#define RT_MSG_DOSERR_80 (RT_MSG_DOSERR + 80)
#define RT_MSG_DOSERR_81 (RT_MSG_DOSERR + 81)
#define RT_MSG_DOSERR_82 (RT_MSG_DOSERR + 82)
#define RT_MSG_DOSERR_83 (RT_MSG_DOSERR + 83)
#define RT_MSG_DOSERR_84 (RT_MSG_DOSERR + 84)
#define RT_MSG_DOSERR_85 (RT_MSG_DOSERR + 85)
#define RT_MSG_DOSERR_86 (RT_MSG_DOSERR + 86)
#define RT_MSG_DOSERR_87 (RT_MSG_DOSERR + 87)
#define RT_MSG_DOSERR_88 (RT_MSG_DOSERR + 88)
#define RT_MSG_DOSERR_89 (RT_MSG_DOSERR + 89)
#define RT_MSG_DOSERR_90 (RT_MSG_DOSERR + 90)
#define RT_MSG_DOSERR_91 (RT_MSG_DOSERR + 91)
#define RT_MSG_DOSERR_92 (RT_MSG_DOSERR + 92)
#define RT_MSG_DOSERR_93 (RT_MSG_DOSERR + 93)
#define RT_MSG_DOSERR_94 (RT_MSG_DOSERR + 94)
#define RT_MSG_DOSERR_95 (RT_MSG_DOSERR + 95)
#define RT_MSG_DOSERR_96 (RT_MSG_DOSERR + 96)
#define RT_MSG_DOSERR_97 (RT_MSG_DOSERR + 97)
#define RT_MSG_DOSERR_98 (RT_MSG_DOSERR + 98)
#define RT_MSG_DOSERR_99 (RT_MSG_DOSERR + 99)
#define RT_MSG_DOSERR_100 (RT_MSG_DOSERR + 100)
#define RT_MSG_DOSERR_101 (RT_MSG_DOSERR + 101)
#define RT_MSG_DOSERR_102 (RT_MSG_DOSERR + 102)
#define RT_MSG_DOSERR_103 (RT_MSG_DOSERR + 103)
#define RT_MSG_DOSERR_104 (RT_MSG_DOSERR + 104)
#define RT_MSG_DOSERR_105 (RT_MSG_DOSERR + 105)
#define RT_MSG_DOSERR_106 (RT_MSG_DOSERR + 106)
#define RT_MSG_DOSERR_107 (RT_MSG_DOSERR + 107)
#define RT_MSG_DOSERR_108 (RT_MSG_DOSERR + 108)
#define RT_MSG_DOSERR_109 (RT_MSG_DOSERR + 109)
#define RT_MSG_DOSERR_110 (RT_MSG_DOSERR + 110)
#define RT_MSG_DOSERR_111 (RT_MSG_DOSERR + 111)
#define RT_MSG_DOSERR_112 (RT_MSG_DOSERR + 112)
#define RT_MSG_DOSERR_113 (RT_MSG_DOSERR + 113)
#define RT_MSG_DOSERR_114 (RT_MSG_DOSERR + 114)
#define RT_MSG_DOSERR_115 (RT_MSG_DOSERR + 115)
#define RT_MSG_DOSERR_116 (RT_MSG_DOSERR + 116)
#define RT_MSG_DOSERR_117 (RT_MSG_DOSERR + 117)
#define RT_MSG_DOSERR_118 (RT_MSG_DOSERR + 118)
#define RT_MSG_DOSERR_119 (RT_MSG_DOSERR + 119)
#define RT_MSG_DOSERR_120 (RT_MSG_DOSERR + 120)
#define RT_MSG_DOSERR_121 (RT_MSG_DOSERR + 121)
#define RT_MSG_DOSERR_122 (RT_MSG_DOSERR + 122)
#define RT_MSG_DOSERR_123 (RT_MSG_DOSERR + 123)
#define RT_MSG_DOSERR_124 (RT_MSG_DOSERR + 124)
#define RT_MSG_DOSERR_125 (RT_MSG_DOSERR + 125)
#define RT_MSG_DOSERR_126 (RT_MSG_DOSERR + 126)
#define RT_MSG_DOSERR_127 (RT_MSG_DOSERR + 127)
#define RT_MSG_DOSERR_128 (RT_MSG_DOSERR + 128)
#define RT_MSG_DOSERR_129 (RT_MSG_DOSERR + 129)
#define RT_MSG_DOSERR_130 (RT_MSG_DOSERR + 130)
#define RT_MSG_DOSERR_131 (RT_MSG_DOSERR + 131)
#define RT_MSG_DOSERR_132 (RT_MSG_DOSERR + 132)
#define RT_MSG_DOSERR_133 (RT_MSG_DOSERR + 133)
#define RT_MSG_DOSERR_134 (RT_MSG_DOSERR + 134)
#define RT_MSG_DOSERR_135 (RT_MSG_DOSERR + 135)
#define RT_MSG_DOSERR_136 (RT_MSG_DOSERR + 136)
#define RT_MSG_DOSERR_137 (RT_MSG_DOSERR + 137)
#define RT_MSG_DOSERR_138 (RT_MSG_DOSERR + 138)
#define RT_MSG_DOSERR_139 (RT_MSG_DOSERR + 139)
#define RT_MSG_DOSERR_140 (RT_MSG_DOSERR + 140)
#define RT_MSG_DOSERR_141 (RT_MSG_DOSERR + 141)
#define RT_MSG_DOSERR_142 (RT_MSG_DOSERR + 142)
#define RT_MSG_DOSERR_143 (RT_MSG_DOSERR + 143)
#define RT_MSG_DOSERR_144 (RT_MSG_DOSERR + 144)
#define RT_MSG_DOSERR_145 (RT_MSG_DOSERR + 145)
#define RT_MSG_DOSERR_146 (RT_MSG_DOSERR + 146)
#define RT_MSG_DOSERR_147 (RT_MSG_DOSERR + 147)
#define RT_MSG_DOSERR_148 (RT_MSG_DOSERR + 148)
#define RT_MSG_DOSERR_149 (RT_MSG_DOSERR + 149)
#define RT_MSG_DOSERR_150 (RT_MSG_DOSERR + 150)
#define RT_MSG_DOSERR_151 (RT_MSG_DOSERR + 151)
#define RT_MSG_DOSERR_152 (RT_MSG_DOSERR + 152)
#define RT_MSG_DOSERR_153 (RT_MSG_DOSERR + 153)
#define RT_MSG_DOSERR_154 (RT_MSG_DOSERR + 154)
#define RT_MSG_DOSERR_155 (RT_MSG_DOSERR + 155)
#define RT_MSG_DOSERR_156 (RT_MSG_DOSERR + 156)
#define RT_MSG_DOSERR_157 (RT_MSG_DOSERR + 157)
#define RT_MSG_DOSERR_158 (RT_MSG_DOSERR + 158)
#define RT_MSG_DOSERR_159 (RT_MSG_DOSERR + 159)
#define RT_MSG_DOSERR_160 (RT_MSG_DOSERR + 160)
#define RT_MSG_DOSERR_161 (RT_MSG_DOSERR + 161)
#define RT_MSG_DOSERR_162 (RT_MSG_DOSERR + 162)
#define RT_MSG_DOSERR_163 (RT_MSG_DOSERR + 163)
#define RT_MSG_DOSERR_164 (RT_MSG_DOSERR + 164)
#define RT_MSG_DOSERR_165 (RT_MSG_DOSERR + 165)
#define RT_MSG_DOSERR_166 (RT_MSG_DOSERR + 166)
#define RT_MSG_DOSERR_167 (RT_MSG_DOSERR + 167)
#define RT_MSG_DOSERR_168 (RT_MSG_DOSERR + 168)
#define RT_MSG_DOSERR_169 (RT_MSG_DOSERR + 169)
#define RT_MSG_DOSERR_170 (RT_MSG_DOSERR + 170)
#define RT_MSG_DOSERR_171 (RT_MSG_DOSERR + 171)
#define RT_MSG_DOSERR_172 (RT_MSG_DOSERR + 172)
#define RT_MSG_DOSERR_173 (RT_MSG_DOSERR + 173)
#define RT_MSG_DOSERR_174 (RT_MSG_DOSERR + 174)
#define RT_MSG_DOSERR_175 (RT_MSG_DOSERR + 175)
#define RT_MSG_DOSERR_176 (RT_MSG_DOSERR + 176)
#define RT_MSG_DOSERR_177 (RT_MSG_DOSERR + 177)
#define RT_MSG_DOSERR_178 (RT_MSG_DOSERR + 178)
#define RT_MSG_DOSERR_179 (RT_MSG_DOSERR + 179)
#define RT_MSG_DOSERR_180 (RT_MSG_DOSERR + 180)
#define RT_MSG_DOSERR_181 (RT_MSG_DOSERR + 181)
#define RT_MSG_DOSERR_182 (RT_MSG_DOSERR + 182)
#define RT_MSG_DOSERR_183 (RT_MSG_DOSERR + 183)
#define RT_MSG_DOSERR_184 (RT_MSG_DOSERR + 184)
#define RT_MSG_DOSERR_185 (RT_MSG_DOSERR + 185)
#define RT_MSG_DOSERR_186 (RT_MSG_DOSERR + 186)
#define RT_MSG_DOSERR_187 (RT_MSG_DOSERR + 187)
#define RT_MSG_DOSERR_188 (RT_MSG_DOSERR + 188)
#define RT_MSG_DOSERR_189 (RT_MSG_DOSERR + 189)
#define RT_MSG_DOSERR_190 (RT_MSG_DOSERR + 190)
#define RT_MSG_DOSERR_191 (RT_MSG_DOSERR + 191)
#define RT_MSG_DOSERR_192 (RT_MSG_DOSERR + 192)
#define RT_MSG_DOSERR_193 (RT_MSG_DOSERR + 193)
#define RT_MSG_DOSERR_194 (RT_MSG_DOSERR + 194)
#define RT_MSG_DOSERR_195 (RT_MSG_DOSERR + 195)
#define RT_MSG_DOSERR_196 (RT_MSG_DOSERR + 196)
#define RT_MSG_DOSERR_197 (RT_MSG_DOSERR + 197)
#define RT_MSG_DOSERR_198 (RT_MSG_DOSERR + 198)
#define RT_MSG_DOSERR_199 (RT_MSG_DOSERR + 199)
#define RT_MSG_DOSERR_200 (RT_MSG_DOSERR + 200)
#define RT_MSG_DOSERR_201 (RT_MSG_DOSERR + 201)
#define RT_MSG_DOSERR_202 (RT_MSG_DOSERR + 202)
#define RT_MSG_DOSERR_203 (RT_MSG_DOSERR + 203)
#define RT_MSG_DOSERR_204 (RT_MSG_DOSERR + 204)
#define RT_MSG_DOSERR_205 (RT_MSG_DOSERR + 205)
#define RT_MSG_DOSERR_206 (RT_MSG_DOSERR + 206)
#define RT_MSG_DOSERR_207 (RT_MSG_DOSERR + 207)
#define RT_MSG_DOSERR_208 (RT_MSG_DOSERR + 208)
#define RT_MSG_DOSERR_209 (RT_MSG_DOSERR + 209)
#define RT_MSG_DOSERR_210 (RT_MSG_DOSERR + 210)
#define RT_MSG_DOSERR_211 (RT_MSG_DOSERR + 211)
#define RT_MSG_DOSERR_212 (RT_MSG_DOSERR + 212)
#define RT_MSG_DOSERR_213 (RT_MSG_DOSERR + 213)
#define RT_MSG_DOSERR_214 (RT_MSG_DOSERR + 214)
#define RT_MSG_DOSERR_215 (RT_MSG_DOSERR + 215)
#define RT_MSG_DOSERR_216 (RT_MSG_DOSERR + 216)
#define RT_MSG_DOSERR_217 (RT_MSG_DOSERR + 217)
#define RT_MSG_DOSERR_218 (RT_MSG_DOSERR + 218)
#define RT_MSG_DOSERR_219 (RT_MSG_DOSERR + 219)
#define RT_MSG_DOSERR_220 (RT_MSG_DOSERR + 220)
#define RT_MSG_DOSERR_221 (RT_MSG_DOSERR + 221)
#define RT_MSG_DOSERR_222 (RT_MSG_DOSERR + 222)
#define RT_MSG_DOSERR_223 (RT_MSG_DOSERR + 223)
#define RT_MSG_DOSERR_224 (RT_MSG_DOSERR + 224)
#define RT_MSG_DOSERR_225 (RT_MSG_DOSERR + 225)
#define RT_MSG_DOSERR_226 (RT_MSG_DOSERR + 226)
#define RT_MSG_DOSERR_227 (RT_MSG_DOSERR + 227)
#define RT_MSG_DOSERR_228 (RT_MSG_DOSERR + 228)
#define RT_MSG_DOSERR_229 (RT_MSG_DOSERR + 229)
#define RT_MSG_DOSERR_230 (RT_MSG_DOSERR + 230)
#define RT_MSG_DOSERR_231 (RT_MSG_DOSERR + 231)
#define RT_MSG_DOSERR_232 (RT_MSG_DOSERR + 232)
#define RT_MSG_DOSERR_233 (RT_MSG_DOSERR + 233)
#define RT_MSG_DOSERR_234 (RT_MSG_DOSERR + 234)
#define RT_MSG_DOSERR_235 (RT_MSG_DOSERR + 235)
#define RT_MSG_DOSERR_236 (RT_MSG_DOSERR + 236)
#define RT_MSG_DOSERR_237 (RT_MSG_DOSERR + 237)
#define RT_MSG_DOSERR_238 (RT_MSG_DOSERR + 238)
#define RT_MSG_DOSERR_239 (RT_MSG_DOSERR + 239)
#define RT_MSG_DOSERR_240 (RT_MSG_DOSERR + 240)
#define RT_MSG_DOSERR_241 (RT_MSG_DOSERR + 241)
#define RT_MSG_DOSERR_242 (RT_MSG_DOSERR + 242)
#define RT_MSG_DOSERR_243 (RT_MSG_DOSERR + 243)
#define RT_MSG_DOSERR_244 (RT_MSG_DOSERR + 244)
#define RT_MSG_DOSERR_245 (RT_MSG_DOSERR + 245)
#define RT_MSG_DOSERR_246 (RT_MSG_DOSERR + 246)
#define RT_MSG_DOSERR_247 (RT_MSG_DOSERR + 247)
#define RT_MSG_DOSERR_248 (RT_MSG_DOSERR + 248)
#define RT_MSG_DOSERR_249 (RT_MSG_DOSERR + 249)
#define RT_MSG_DOSERR_250 (RT_MSG_DOSERR + 250)
#define RT_MSG_DOSERR_251 (RT_MSG_DOSERR + 251)
#define RT_MSG_DOSERR_252 (RT_MSG_DOSERR + 252)
#define RT_MSG_DOSERR_253 (RT_MSG_DOSERR + 253)
#define RT_MSG_DOSERR_254 (RT_MSG_DOSERR + 254)
#define RT_MSG_DOSERR_255 (RT_MSG_DOSERR + 255)
#define RT_MSG_DOSERR_256 (RT_MSG_DOSERR + 256)
#define RT_MSG_DOSERR_257 (RT_MSG_DOSERR + 257)
#define RT_MSG_DOSERR_258 (RT_MSG_DOSERR + 258)
#define RT_MSG_DOSERR_FFFF (RT_MSG_DOSERR + 259)
#define RT_MSG_DOSERR_UNKNOW (RT_MSG_DOSERR + 260)
#define __CAVOSTR_SYSLIB_FIRST_STRING 5000
#define __CAVOSTR_SYSLIB_LAST_STRING 5099
#define __CAVOSTR_SYSLIB_ARG (__CAVOSTR_SYSLIB_FIRST_STRING+ 2)
#define __CAVOSTR_SYSLIB_ARG_ERROR (__CAVOSTR_SYSLIB_FIRST_STRING+ 3)
#define __CAVOSTR_SYSLIB_ARGNUM (__CAVOSTR_SYSLIB_FIRST_STRING+ 4)
#define __CAVOSTR_SYSLIB_ARGS (__CAVOSTR_SYSLIB_FIRST_STRING+ 5)
#define __CAVOSTR_SYSLIB_ARGTYPE (__CAVOSTR_SYSLIB_FIRST_STRING+ 6)
#define __CAVOSTR_SYSLIB_ARGTYPE_REQ (__CAVOSTR_SYSLIB_FIRST_STRING+ 7)
#define __CAVOSTR_SYSLIB_BADTRANSLATIONARRAY (__CAVOSTR_SYSLIB_FIRST_STRING+ 1)
#define __CAVOSTR_SYSLIB_CALLED_FROM (__CAVOSTR_SYSLIB_FIRST_STRING+ 8)
#define __CAVOSTR_SYSLIB_CHOICE (__CAVOSTR_SYSLIB_FIRST_STRING+ 9)
#define __CAVOSTR_SYSLIB_CMD_LINE (__CAVOSTR_SYSLIB_FIRST_STRING+10)
#define __CAVOSTR_SYSLIB_CONVERSION (__CAVOSTR_SYSLIB_FIRST_STRING+11)
#define __CAVOSTR_SYSLIB_CURDIR (__CAVOSTR_SYSLIB_FIRST_STRING+12)
#define __CAVOSTR_SYSLIB_DANGER (__CAVOSTR_SYSLIB_FIRST_STRING+13)
#define __CAVOSTR_SYSLIB_DISK (__CAVOSTR_SYSLIB_FIRST_STRING+14)
#define __CAVOSTR_SYSLIB_DISK_FREE (__CAVOSTR_SYSLIB_FIRST_STRING+15)
#define __CAVOSTR_SYSLIB_DOS_ERROR (__CAVOSTR_SYSLIB_FIRST_STRING+16)
#define __CAVOSTR_SYSLIB_ENTITY (__CAVOSTR_SYSLIB_FIRST_STRING+17)
#define __CAVOSTR_SYSLIB_ERR_IN_ERR (__CAVOSTR_SYSLIB_FIRST_STRING+18)
#define __CAVOSTR_SYSLIB_ERROR (__CAVOSTR_SYSLIB_FIRST_STRING+19)
#define __CAVOSTR_SYSLIB_FILE (__CAVOSTR_SYSLIB_FIRST_STRING+20)
#define __CAVOSTR_SYSLIB_FILE_HANDLE (__CAVOSTR_SYSLIB_FIRST_STRING+21)
#define __CAVOSTR_SYSLIB_FUNCPTR (__CAVOSTR_SYSLIB_FIRST_STRING+22)
#define __CAVOSTR_SYSLIB_FUNCTION (__CAVOSTR_SYSLIB_FIRST_STRING+23)
#define __CAVOSTR_SYSLIB_HANDLE (__CAVOSTR_SYSLIB_FIRST_STRING+24)
#define __CAVOSTR_SYSLIB_HANDLE_CUR (__CAVOSTR_SYSLIB_FIRST_STRING+25)
#define __CAVOSTR_SYSLIB_HANDLE_END (__CAVOSTR_SYSLIB_FIRST_STRING+26)
#define __CAVOSTR_SYSLIB_IVARS (__CAVOSTR_SYSLIB_FIRST_STRING+27)
#define __CAVOSTR_SYSLIB_LINE (__CAVOSTR_SYSLIB_FIRST_STRING+28)
#define __CAVOSTR_SYSLIB_MAX (__CAVOSTR_SYSLIB_FIRST_STRING+29)
#define __CAVOSTR_SYSLIB_MODULE (__CAVOSTR_SYSLIB_FIRST_STRING+30)
#define __CAVOSTR_SYSLIB_OBJECT (__CAVOSTR_SYSLIB_FIRST_STRING+31)
#define __CAVOSTR_SYSLIB_OPERATION (__CAVOSTR_SYSLIB_FIRST_STRING+32)
#define __CAVOSTR_SYSLIB_SUBCODE (__CAVOSTR_SYSLIB_FIRST_STRING+33)
#define __CAVOSTR_SYSLIB_SUBST_TYPE (__CAVOSTR_SYSLIB_FIRST_STRING+34)
#define __CAVOSTR_SYSLIB_SUBSYSTEM (__CAVOSTR_SYSLIB_FIRST_STRING+35)
#define __CAVOSTR_SYSLIB_TO (__CAVOSTR_SYSLIB_FIRST_STRING+36)
#define __CAVOSTR_SYSLIB_TRIES (__CAVOSTR_SYSLIB_FIRST_STRING+37)
#define __CAVOSTR_SYSLIB_WARNING (__CAVOSTR_SYSLIB_FIRST_STRING+38)
#define __CAVOSTR_SYSLIB_OLEBASE (__CAVOSTR_SYSLIB_FIRST_STRING+39)
#define __CAVOSTR_SYSLIB_CONVERSION_CALLED_FROM (__CAVOSTR_SYSLIB_FIRST_STRING+40)
#define __CAVOSTR_SYSLIB_CONVERSION_TO (__CAVOSTR_SYSLIB_FIRST_STRING+41)
#define __CAVOSTR_SYSLIB_CONVERSION_TO_CALLED_FROM (__CAVOSTR_SYSLIB_FIRST_STRING+42)
#define __CAVOSTR_SYSLIB_FUNCTION_CALLED_FROM (__CAVOSTR_SYSLIB_FIRST_STRING+43)
#define __CAVOSTR_SYSLIB_NOMEM (__CAVOSTR_SYSLIB_FIRST_STRING+44)
#define __CAVOSTR_SYSLIB_INCTYPES (__CAVOSTR_SYSLIB_FIRST_STRING+45)
#define __CAVOSTR_SYSCLASS_FIRST_STRING 5100
#define __CAVOSTR_SYSCLASS_LAST_STRING 5199
#define __CAVOSTR_SYSCLASS_BADDESCRIPTION (__CAVOSTR_SYSCLASS_FIRST_STRING+3)
#define __CAVOSTR_SYSCLASS_BADCAPTION (__CAVOSTR_SYSCLASS_FIRST_STRING+2)
#define __CAVOSTR_SYSCLASS_BADERROROBJECT (__CAVOSTR_SYSCLASS_FIRST_STRING+1)
#define __CAVOSTR_SYSCLASS_BADHELPCONTEXT (__CAVOSTR_SYSCLASS_FIRST_STRING+4)
#define __CAVOSTR_SYSCLASS_BADNAME (__CAVOSTR_SYSCLASS_FIRST_STRING+5)
#define __CAVOSTR_DBFCLASS_FIRST_STRING 5200
#define __CAVOSTR_DBFCLASS_LAST_STRING 5299
#define __CAVOSTR_DBFCLASS_SELECTIVEVALUE (__CAVOSTR_DBFCLASS_FIRST_STRING+32)
#define __CAVOSTR_DBFCLASS_ALIAS (__CAVOSTR_DBFCLASS_FIRST_STRING+1)
#define __CAVOSTR_DBFCLASS_BADCB (__CAVOSTR_DBFCLASS_FIRST_STRING+38)
#define __CAVOSTR_DBFCLASS_BADCHILD (__CAVOSTR_DBFCLASS_FIRST_STRING+2)
#define __CAVOSTR_DBFCLASS_BADCONCURRENCYASSIGN (__CAVOSTR_DBFCLASS_FIRST_STRING+35)
#define __CAVOSTR_DBFCLASS_BADDECIMALS (__CAVOSTR_DBFCLASS_FIRST_STRING+39)
#define __CAVOSTR_DBFCLASS_BADDRIVE (__CAVOSTR_DBFCLASS_FIRST_STRING+40)
#define __CAVOSTR_DBFCLASS_BADEXPRESSION (__CAVOSTR_DBFCLASS_FIRST_STRING+3)
#define __CAVOSTR_DBFCLASS_BADEXTENSION (__CAVOSTR_DBFCLASS_FIRST_STRING+41)
#define __CAVOSTR_DBFCLASS_BADFIELDMATCH (__CAVOSTR_DBFCLASS_FIRST_STRING+4)
#define __CAVOSTR_DBFCLASS_BADFIELDPOSITION (__CAVOSTR_DBFCLASS_FIRST_STRING+36)
#define __CAVOSTR_DBFCLASS_BADFILENAME (__CAVOSTR_DBFCLASS_FIRST_STRING+5)
#define __CAVOSTR_DBFCLASS_BADFILTERBLOCK (__CAVOSTR_DBFCLASS_FIRST_STRING+6)
#define __CAVOSTR_DBFCLASS_BADFS (__CAVOSTR_DBFCLASS_FIRST_STRING+33)
#define __CAVOSTR_DBFCLASS_BADHL (__CAVOSTR_DBFCLASS_FIRST_STRING+42)
#define __CAVOSTR_DBFCLASS_BADHLNAME (__CAVOSTR_DBFCLASS_FIRST_STRING+34)
#define __CAVOSTR_DBFCLASS_BADLENGTH (__CAVOSTR_DBFCLASS_FIRST_STRING+43)
#define __CAVOSTR_DBFCLASS_BADLREQ (__CAVOSTR_DBFCLASS_FIRST_STRING+44)
#define __CAVOSTR_DBFCLASS_BADNAME (__CAVOSTR_DBFCLASS_FIRST_STRING+45)
#define __CAVOSTR_DBFCLASS_BADNEXT (__CAVOSTR_DBFCLASS_FIRST_STRING+7)
#define __CAVOSTR_DBFCLASS_BADNEXT_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+8)
#define __CAVOSTR_DBFCLASS_BADPATH (__CAVOSTR_DBFCLASS_FIRST_STRING+46)
#define __CAVOSTR_DBFCLASS_BADREADONLYMODE (__CAVOSTR_DBFCLASS_FIRST_STRING+9)
#define __CAVOSTR_DBFCLASS_BADSHAREMODE (__CAVOSTR_DBFCLASS_FIRST_STRING+10)
#define __CAVOSTR_DBFCLASS_BADSI (__CAVOSTR_DBFCLASS_FIRST_STRING+47)
#define __CAVOSTR_DBFCLASS_BADSTRING (__CAVOSTR_DBFCLASS_FIRST_STRING+48)
#define __CAVOSTR_DBFCLASS_BADTRANSLATIONARRAY (__CAVOSTR_DBFCLASS_FIRST_STRING+37)
#define __CAVOSTR_DBFCLASS_BADTYPE (__CAVOSTR_DBFCLASS_FIRST_STRING+49)
#define __CAVOSTR_DBFCLASS_BADTYPE2 (__CAVOSTR_DBFCLASS_FIRST_STRING+50)
#define __CAVOSTR_DBFCLASS_FIELDSPEC (__CAVOSTR_DBFCLASS_FIRST_STRING+11)
#define __CAVOSTR_DBFCLASS_INVALIDLENGTH (__CAVOSTR_DBFCLASS_FIRST_STRING+51)
#define __CAVOSTR_DBFCLASS_INVALIDMAX (__CAVOSTR_DBFCLASS_FIRST_STRING+52)
#define __CAVOSTR_DBFCLASS_INVALIDMIN (__CAVOSTR_DBFCLASS_FIRST_STRING+53)
#define __CAVOSTR_DBFCLASS_INVALIDMINLENGTH (__CAVOSTR_DBFCLASS_FIRST_STRING+54)
#define __CAVOSTR_DBFCLASS_INVALIDRANGE (__CAVOSTR_DBFCLASS_FIRST_STRING+55)
#define __CAVOSTR_DBFCLASS_INVALIDTYPE (__CAVOSTR_DBFCLASS_FIRST_STRING+57)
#define __CAVOSTR_DBFCLASS_INVALIDVALUE (__CAVOSTR_DBFCLASS_FIRST_STRING+58)
#define __CAVOSTR_DBFCLASS_LOCKFAILED (__CAVOSTR_DBFCLASS_FIRST_STRING+12)
#define __CAVOSTR_DBFCLASS_LOCKFAILED_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+13)
#define __CAVOSTR_DBFCLASS_MISMATCH (__CAVOSTR_DBFCLASS_FIRST_STRING+14)
#define __CAVOSTR_DBFCLASS_NODATAFIELDSEXIST (__CAVOSTR_DBFCLASS_FIRST_STRING+15)
#define __CAVOSTR_DBFCLASS_NOFIELDS (__CAVOSTR_DBFCLASS_FIRST_STRING+16)
#define __CAVOSTR_DBFCLASS_NOFILENAME (__CAVOSTR_DBFCLASS_FIRST_STRING+17)
#define __CAVOSTR_DBFCLASS_NOGOTOP (__CAVOSTR_DBFCLASS_FIRST_STRING+18)
#define __CAVOSTR_DBFCLASS_NOGOTOP_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+19)
#define __CAVOSTR_DBFCLASS_NOSEEK (__CAVOSTR_DBFCLASS_FIRST_STRING+20)
#define __CAVOSTR_DBFCLASS_NOSELECTIONACTIVE (__CAVOSTR_DBFCLASS_FIRST_STRING+21)
#define __CAVOSTR_DBFCLASS_NOTABLE (__CAVOSTR_DBFCLASS_FIRST_STRING+22)
#define __CAVOSTR_DBFCLASS_NOTABLE_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+23)
#define __CAVOSTR_DBFCLASS_NOTABLE2 (__CAVOSTR_DBFCLASS_FIRST_STRING+24)
#define __CAVOSTR_DBFCLASS_RECORDCHANGED (__CAVOSTR_DBFCLASS_FIRST_STRING+25)
#define __CAVOSTR_DBFCLASS_RECORDCHANGED_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+26)
#define __CAVOSTR_DBFCLASS_REQUIRED (__CAVOSTR_DBFCLASS_FIRST_STRING+59)
#define __CAVOSTR_DBFCLASS_SELECTIVENOTFOUND (__CAVOSTR_DBFCLASS_FIRST_STRING+30)
#define __CAVOSTR_DBFCLASS_SELECTIVESEEK (__CAVOSTR_DBFCLASS_FIRST_STRING+31)
#define __CAVOSTR_DBFCLASS_INTENTTOMOVE (__CAVOSTR_DBFCLASS_FIRST_STRING+60)
#define __CAVOSTR_DBFCLASS_INTENTTOMOVE_CAPTION (__CAVOSTR_DBFCLASS_FIRST_STRING+61)
#define __CAVOSTR_DBFCLASS_BADPARENT (__CAVOSTR_DBFCLASS_FIRST_STRING+62)
#define __CAVOSTR_DBFCLASS_INVALIDINDEX (__CAVOSTR_DBFCLASS_FIRST_STRING+63)
#define __CAVOSTR_DBFCLASS_KEYVALUE (__CAVOSTR_DBFCLASS_FIRST_STRING+64)
#define __CAVOSTR_DBFCLASS_INVALIDORDER (__CAVOSTR_DBFCLASS_FIRST_STRING+65)
#define __CAVOSTR_DBFCLASS_NOFIELDMATCH (__CAVOSTR_DBFCLASS_FIRST_STRING+66)
#define __CAVOSTR_DBFCLASS_BADALIAS (__CAVOSTR_DBFCLASS_FIRST_STRING+67)
#define __CAVOSTR_DBFCLASS_BADERROROBJECT (__CAVOSTR_DBFCLASS_FIRST_STRING+68)
#define OLEAUTO_ERROR_FIRST 5300
#define OLEAUTO_ERROR_LAST (OLEAUTO_ERROR_FIRST + 100)
#define OLEAUTO_ERROR_SUBSYSTEM (OLEAUTO_ERROR_FIRST + 0)
#define OLEAUTO_ERROR_MSG_NO_GET_PROPERTY (OLEAUTO_ERROR_FIRST + 1)
#define OLEAUTO_ERROR_MSG_NO_SET_PROPERTY (OLEAUTO_ERROR_FIRST + 2)
#define OLEAUTO_ERROR_MSG_UNKNOWN_ERROR (OLEAUTO_ERROR_FIRST + 3)
#define OLEAUTO_ERROR_MSG_NO_MEMORY (OLEAUTO_ERROR_FIRST + 4)
#define OLEAUTO_ERROR_MSG_CONVERTERR (OLEAUTO_ERROR_FIRST + 5)
#define OLEAUTO_ERROR_EXP_NO_DESC (OLEAUTO_ERROR_FIRST + 6)
#define OLEAUTO_ERROR_MSG_GET_PROPERTY_FAILED (OLEAUTO_ERROR_FIRST + 7)
#define OLEAUTO_ERROR_MSG_SET_PROPERTY_FAILED (OLEAUTO_ERROR_FIRST + 8)
#define OLEAUTO_ERROR_MSG_NO_METHOD (OLEAUTO_ERROR_FIRST + 9)
#define OLEAUTO_ERROR_MSG_METHOD_FAILED (OLEAUTO_ERROR_FIRST + 10)
#define OLEAUTO_ERROR_MSG_PARAM_MISSING (OLEAUTO_ERROR_FIRST + 11)
#define OLEAUTO_ERROR_MSG_NAMED_ARG (OLEAUTO_ERROR_FIRST + 12)
#define OLEAUTO_ERROR_MSG_INIT_FAILED (OLEAUTO_ERROR_FIRST + 13)
#define OLEAUTO_ERROR_MSG_NAMED_ARG_LAST (OLEAUTO_ERROR_FIRST + 14)
#define OLEAUTO_ERROR_MSG_NAMED_ARG_NOTSUPP (OLEAUTO_ERROR_FIRST + 15)
#define OLEAUTO_ERROR_MSG_VARIANT_ARGS (OLEAUTO_ERROR_FIRST + 16)
#define OLEAUTO_ERROR_NO_IDISPATCH_INTERFACE (OLEAUTO_ERROR_FIRST + 17)
#define OLEAUTO_ERROR_NO_ITYPELIB_INTERFACE (OLEAUTO_ERROR_FIRST + 18)
#define IDS_OLERUNTIME (OLEAUTO_ERROR_FIRST + 50)
#define IDS_NOAPPDOCFILE (OLEAUTO_ERROR_FIRST + 51)
#define IDS_NOINSERT (OLEAUTO_ERROR_FIRST + 52)
#define IDS_CREATEFAILED (OLEAUTO_ERROR_FIRST + 53)
#define __CAVOSTR_GUICLASS_FIRST_STRING 5400
#define __CAVOSTR_GUICLASS_LAST_STRING 5499
#define __CAVOSTR_GUICLASS_ASSERTFAILED (__CAVOSTR_GUICLASS_FIRST_STRING+ 1)
#define __CAVOSTR_GUICLASS_ASSERTIONFAILED (__CAVOSTR_GUICLASS_FIRST_STRING+ 2)
#define __CAVOSTR_GUICLASS_ATTEMPTREPORTS (__CAVOSTR_GUICLASS_FIRST_STRING+ 3)
#define __CAVOSTR_GUICLASS_CAPTIONINVALID (__CAVOSTR_GUICLASS_FIRST_STRING+ 7)
#define __CAVOSTR_GUICLASS_CHANGINGVIEW (__CAVOSTR_GUICLASS_FIRST_STRING+ 8)
#define __CAVOSTR_GUICLASS_CHGDISCARD (__CAVOSTR_GUICLASS_FIRST_STRING+ 9)
#define __CAVOSTR_GUICLASS_CLOSINGCHANGES (__CAVOSTR_GUICLASS_FIRST_STRING+10)
#define __CAVOSTR_GUICLASS_CLOSINGINVCHANGES (__CAVOSTR_GUICLASS_FIRST_STRING+11)
#define __CAVOSTR_GUICLASS_CVIDINVALID (__CAVOSTR_GUICLASS_FIRST_STRING+13)
#define __CAVOSTR_GUICLASS_DATAWINDOW (__CAVOSTR_GUICLASS_FIRST_STRING+14)
#define __CAVOSTR_GUICLASS_DBROWSEROBJEDT (__CAVOSTR_GUICLASS_FIRST_STRING+15)
#define __CAVOSTR_GUICLASS_DELETEDRECORD (__CAVOSTR_GUICLASS_FIRST_STRING+16)
#define __CAVOSTR_GUICLASS_DELETEFAILED (__CAVOSTR_GUICLASS_FIRST_STRING+17)
#define __CAVOSTR_GUICLASS_DELETEFAILEDMSG (__CAVOSTR_GUICLASS_FIRST_STRING+18)
#define __CAVOSTR_GUICLASS_DWUNTITLED (__CAVOSTR_GUICLASS_FIRST_STRING+19)
#define __CAVOSTR_GUICLASS_ERROR (__CAVOSTR_GUICLASS_FIRST_STRING+20)
#define __CAVOSTR_GUICLASS_INTERFACEERROR (__CAVOSTR_GUICLASS_FIRST_STRING+22)
#define __CAVOSTR_GUICLASS_INVALIDARG (__CAVOSTR_GUICLASS_FIRST_STRING+23)
#define __CAVOSTR_GUICLASS_INVALIDCAT (__CAVOSTR_GUICLASS_FIRST_STRING+24)
#define __CAVOSTR_GUICLASS_INVALIDRPC (__CAVOSTR_GUICLASS_FIRST_STRING+25)
#define __CAVOSTR_GUICLASS_INVALIDVIEW (__CAVOSTR_GUICLASS_FIRST_STRING+26)
#define __CAVOSTR_GUICLASS_INVARGUMENT (__CAVOSTR_GUICLASS_FIRST_STRING+27)
#define __CAVOSTR_GUICLASS_INVMETHODARG (__CAVOSTR_GUICLASS_FIRST_STRING+28)
#define __CAVOSTR_GUICLASS_NOPROMPT (__CAVOSTR_GUICLASS_FIRST_STRING+29)
#define __CAVOSTR_GUICLASS_NOTFOUND (__CAVOSTR_GUICLASS_FIRST_STRING+30)
#define __CAVOSTR_GUICLASS_OWNERINVALID (__CAVOSTR_GUICLASS_FIRST_STRING+31)
#define __CAVOSTR_GUICLASS_PARMINVALID (__CAVOSTR_GUICLASS_FIRST_STRING+32)
#define __CAVOSTR_GUICLASS_SHOULDAPP (__CAVOSTR_GUICLASS_FIRST_STRING+33)
#define __CAVOSTR_GUICLASS_TYPEERROR (__CAVOSTR_GUICLASS_FIRST_STRING+34)
#define __CAVOSTR_GUICLASS_UNKNOWN (__CAVOSTR_GUICLASS_FIRST_STRING+36)
#define __CAVOSTR_GUICLASS_UNKNOWNPARM (__CAVOSTR_GUICLASS_FIRST_STRING+37)
#define __CAVOSTR_GUICLASS_UNKNOWNSTATUS (__CAVOSTR_GUICLASS_FIRST_STRING+38)
#define __CAVOSTR_GUICLASS_UNKNOWNSTATUSMSG (__CAVOSTR_GUICLASS_FIRST_STRING+39)
#define __CAVOSTR_GUICLASS_WARNING (__CAVOSTR_GUICLASS_FIRST_STRING+40)
#define __CAVOSTR_GUICLASS_WARNING2 (__CAVOSTR_GUICLASS_FIRST_STRING+41)
#define __CAVOSTR_GUICLASS_WARNING3 (__CAVOSTR_GUICLASS_FIRST_STRING+42)
#define __CAVOSTR_GUICLASS_YOUHAVECLOSED (__CAVOSTR_GUICLASS_FIRST_STRING+43)
#define __CAVOSTR_GUICLASS_ERROR2 (__CAVOSTR_GUICLASS_FIRST_STRING+44)
#define __CAVOSTR_GUICLASS_INFO (__CAVOSTR_GUICLASS_FIRST_STRING+45)
#define __CAVOSTR_GUICLASS_DSNOTOPEN (__CAVOSTR_GUICLASS_FIRST_STRING+46)
#define __WCSFirst 4000
#define __WCSLibraryName (__WCSFirst + 1)
#define __WCSInterfaceError (__WCSFirst + 2)
#define __WCSTypeError (__WCSFirst + 3)
#define __WCSLoadLibraryError (__WCSFirst + 4)
#define __WCSError (__WCSFirst + 5)
#define __WCSAreaIndex (__WCSFirst + 6)
#define __WCSAreaIndexLast (__WCSFirst + 30)
#define __WCSUnknown (__WCSFirst + 31)
#define __WCSWarning (__WCSFirst + 32)
#define __WCSChgDiscard (__WCSFirst + 33)
#define __WCSDataWindow (__WCSFirst + 34)
#define __WCSDWUntitled (__WCSFirst + 35)
#define __WCSUnknownStatus (__WCSFirst + 36)
#define __WCSUnknownStatusMSG (__WCSFirst + 37)
#define __WCSError2 (__WCSFirst + 38)
#define __WCSDSNotOpen (__WCSFirst + 39)
#define __WCSChangingView (__WCSFirst + 41)
#define __WCSDeletedRecord (__WCSFirst + 43)
#define __WCSIpcServerNotFound (__WCSFirst + 44)
#define __WCSIpcTopicNotFound (__WCSFirst + 45)
#define __WCSIpcItemNotFound (__WCSFirst + 46)
#define __WCSIpcOutOfMemory (__WCSFirst + 47)
#define __WCSDeleteFailed (__WCSFirst + 40)
#define __WCSDeleteFailedMSG (__WCSFirst + 42)
#define __WCSAllFiles (__WCSFirst + 48)
#define __WCSPrinterNoDiskSpace (__WCSFirst + 49)
#define __WCSDataDialog (__WCSFirst + 50)
#define __WCSDBrowserObject (__WCSFirst + 51)
#define __WCSCreateCtlFailed (__WCSFirst + 52)
#define __WCSCreateDlgFailed (__WCSFirst + 53)
#define __WCSHostVOApp (__WCSFirst + 54)
#define __WCSHostDataBrowser (__WCSFirst + 55)
#define __WCSHostDataWindow (__WCSFirst + 56)
#define __WCSPictureYN (__WCSFirst + 57)
#define __WCSPictureTFYN (__WCSFirst + 58)
#define __WCSNoOLESupport (__WCSFirst + 59)
#define __WCSTextBox (__WCSFirst + 60)
#define __WCSInfoBox (__WCSFirst + 61)
#define __WCSCAPaintLoadFailed (__WCSFirst + 62)
#define __WCSCNoAutomation (__WCSFirst + 63)
#define __WCToolBarOffset (__WCSFirst + 64)
#define __WCSLast 4999
#define __WCToolTipOffset (__WCToolBarOffset + 134)
#define __CAVOSTR_REPORTCLASS_FIRST_STRING 5500
#define __CAVOSTR_REPORTCLASS_LAST_STRING 5599
#define __CAVOSTR_REPORTCLASS_CLOSEDREPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 2)
#define __CAVOSTR_REPORTCLASS_COMMANDERROR1 (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 3)
#define __CAVOSTR_REPORTCLASS_COMMANDERROR2 (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 4)
#define __CAVOSTR_REPORTCLASS_COMPLETEDREPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 5)
#define __CAVOSTR_REPORTCLASS_DETECTEDERRORS (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 6)
#define __CAVOSTR_REPORTCLASS_OPENEDREPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 7)
#define __CAVOSTR_REPORTCLASS_SAVEDREPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 8)
#define __CAVOSTR_REPORTCLASS_SAVETOFILEINFO1 (__CAVOSTR_REPORTCLASS_FIRST_STRING+ 9)
#define __CAVOSTR_REPORTCLASS_SAVETOFILEINFO2 (__CAVOSTR_REPORTCLASS_FIRST_STRING+10)
#define __CAVOSTR_REPORTCLASS_THEREPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+11)
#define __CAVOSTR_REPORTCLASS_TOCLOSEFILE (__CAVOSTR_REPORTCLASS_FIRST_STRING+12)
#define __CAVOSTR_REPORTCLASS_SYNCHRONOUS (__CAVOSTR_REPORTCLASS_FIRST_STRING+13)
#define __CAVOSTR_REPORTCLASS_ASYNCHRONOUS (__CAVOSTR_REPORTCLASS_FIRST_STRING+14)
#define __CAVOSTR_REPORTCLASS_DDE_PENDING (__CAVOSTR_REPORTCLASS_FIRST_STRING+15)
#define __CAVOSTR_REPORTCLASS_REPORTS_OPEN (__CAVOSTR_REPORTCLASS_FIRST_STRING+16)
#define __CAVOSTR_REPORTCLASS_REPORT (__CAVOSTR_REPORTCLASS_FIRST_STRING+17)
#define __CAVOSTR_REPORTCLASS_ISCLOSED (__CAVOSTR_REPORTCLASS_FIRST_STRING+18)
#define __CAVOSTR_REPORTCLASS_ABOUTTITLE (__CAVOSTR_REPORTCLASS_FIRST_STRING+19)
#define __CAVOSTR_REPORTCLASS_ABOUTBODY (__CAVOSTR_REPORTCLASS_FIRST_STRING+20)
#define __CAVOSTR_REPORTCLASS_PARAMERROR (__CAVOSTR_REPORTCLASS_FIRST_STRING+21)
#define __CAVOSTR_SQLCLASS_FIRST_STRING 5600
#define __CAVOSTR_SQLCLASS_LAST_STRING 5699
#define __CAVOSTR_SQLCLASS_SUBSYS (__CAVOSTR_SQLCLASS_FIRST_STRING+ 1)
#define __CAVOSTR_SQLCLASS__ENV_ALLOC (__CAVOSTR_SQLCLASS_FIRST_STRING+ 2)
#define __CAVOSTR_SQLCLASS__ENV_FREE (__CAVOSTR_SQLCLASS_FIRST_STRING+ 3)
#define __CAVOSTR_SQLCLASS__CON_ALLOC (__CAVOSTR_SQLCLASS_FIRST_STRING+ 4)
#define __CAVOSTR_SQLCLASS__CON_FREE (__CAVOSTR_SQLCLASS_FIRST_STRING+ 5)
#define __CAVOSTR_SQLCLASS__CONNECTED (__CAVOSTR_SQLCLASS_FIRST_STRING+ 6)
#define __CAVOSTR_SQLCLASS__NOT_CONN (__CAVOSTR_SQLCLASS_FIRST_STRING+ 7)
#define __CAVOSTR_SQLCLASS__CANCELLED (__CAVOSTR_SQLCLASS_FIRST_STRING+ 9)
#define __CAVOSTR_SQLCLASS__ODBC_VO (__CAVOSTR_SQLCLASS_FIRST_STRING+10)
#define __CAVOSTR_SQLCLASS__GENERAL_ERR (__CAVOSTR_SQLCLASS_FIRST_STRING+11)
#define __CAVOSTR_SQLCLASS__STMT_NOT_ALLOC (__CAVOSTR_SQLCLASS_FIRST_STRING+12)
#define __CAVOSTR_SQLCLASS__STMT_PREP (__CAVOSTR_SQLCLASS_FIRST_STRING+13)
#define __CAVOSTR_SQLCLASS__NO_STMT (__CAVOSTR_SQLCLASS_FIRST_STRING+14)
#define __CAVOSTR_SQLCLASS__STMT_ALLOC (__CAVOSTR_SQLCLASS_FIRST_STRING+15)
#define __CAVOSTR_SQLCLASS__FUNCSEQ_ERR (__CAVOSTR_SQLCLASS_FIRST_STRING+16)
#define __CAVOSTR_SQLCLASS__PARM_TYPE (__CAVOSTR_SQLCLASS_FIRST_STRING+17)
#define __CAVOSTR_SQLCLASS__MEM_ALLOC (__CAVOSTR_SQLCLASS_FIRST_STRING+18)
#define __CAVOSTR_SQLCLASS__BADCOL (__CAVOSTR_SQLCLASS_FIRST_STRING+19)
#define __CAVOSTR_SQLCLASS__BADFLD (__CAVOSTR_SQLCLASS_FIRST_STRING+20)
#define __CAVOSTR_SQLCLASS__BADPAR (__CAVOSTR_SQLCLASS_FIRST_STRING+21)
#define __CAVOSTR_SQLCLASS__BADRECNO (__CAVOSTR_SQLCLASS_FIRST_STRING+22)
#define __CAVOSTR_SQLCLASS__BACKWARDS (__CAVOSTR_SQLCLASS_FIRST_STRING+23)
#define __CAVOSTR_SQLCLASS__BOF (__CAVOSTR_SQLCLASS_FIRST_STRING+24)
#define __CAVOSTR_SQLCLASS__EOF (__CAVOSTR_SQLCLASS_FIRST_STRING+25)
#define __CAVOSTR_SQLCLASS__NOFLDS (__CAVOSTR_SQLCLASS_FIRST_STRING+26)
#define __CAVOSTR_SQLCLASS__NO_KEY (__CAVOSTR_SQLCLASS_FIRST_STRING+27)
#define __CAVOSTR_SQLCLASS__NO_ROW (__CAVOSTR_SQLCLASS_FIRST_STRING+28)
#define __CAVOSTR_SQLCLASS__NO_INS (__CAVOSTR_SQLCLASS_FIRST_STRING+29)
#define __CAVOSTR_SQLCLASS__INV_OP (__CAVOSTR_SQLCLASS_FIRST_STRING+30)
#define __CAVOSTR_SQLCLASS__NO_CSR (__CAVOSTR_SQLCLASS_FIRST_STRING+31)
#define __CAVOSTR_SQLCLASS__BADVALID (__CAVOSTR_SQLCLASS_FIRST_STRING+32)
#define __CAVOSTR_SQLCLASS__EMPTY (__CAVOSTR_SQLCLASS_FIRST_STRING+33)
#define __CAVOSTR_SQLCLASS__UPDATE_COL (__CAVOSTR_SQLCLASS_FIRST_STRING+34)
#define __CAVOSTR_SQLCLASS__NODATAFIELDSEXIST (__CAVOSTR_SQLCLASS_FIRST_STRING+35)
#define __CAVOSTR_SQLCLASS__BADFIELDPOSITION (__CAVOSTR_SQLCLASS_FIRST_STRING+36)
#define __CAVOSTR_SQLCLASS__INVALIDCOLATT (__CAVOSTR_SQLCLASS_FIRST_STRING+37)
#define TERMINAL_FIRST 5700
#define TERMINAL_LAST 5799
#define TMSG_YN (TERMINAL_FIRST + 1)
#define TMSG_ALERTDEFAULT (TERMINAL_FIRST + 2)
#define TMSG_NOTERMWIN (TERMINAL_FIRST + 3)
#define TMSG_FNTCHNG (TERMINAL_FIRST + 4)
#define TMSG_SHADE (TERMINAL_FIRST + 5)
#define TMSG_MARK (TERMINAL_FIRST + 6)
#define TMSG_SCREEN2FILE (TERMINAL_FIRST + 7)
#define TMSG_MEMRECOUR (TERMINAL_FIRST + 8)
#define TMSG_DYNCHECKERR (TERMINAL_FIRST + 9)
#define TMSG_HNDLINE (TERMINAL_FIRST + 10)
#define TMSG_HNDENTITY (TERMINAL_FIRST + 11)
#define TMSG_HNDCONTENTS (TERMINAL_FIRST + 12)
#define TMSG_HNDVAR (TERMINAL_FIRST + 13)
#define TMSG_NOCHANGE (TERMINAL_FIRST + 14)
#define TMSG_FONTCHGERR (TERMINAL_FIRST + 15)
#define TMSG_MUSTSELECT (TERMINAL_FIRST + 16)
#define TMSG_NODEVSEL (TERMINAL_FIRST + 17)
#define TMSG_NOLINK (TERMINAL_FIRST + 18)
#define TMSG_PRNSETUP (TERMINAL_FIRST + 19)
#define TMSG_PAGENO (TERMINAL_FIRST + 20)
#define TMSG_PRESSANYKEY (TERMINAL_FIRST + 21)
#define TMSG_APPENDSCREEN (TERMINAL_FIRST + 22)
#define TMSG_APPENDALL (TERMINAL_FIRST + 23)
#define TMSG_LOCKEDFONT (TERMINAL_FIRST + 24)
#define TMSG_NOACCELERATORS (TERMINAL_FIRST + 25)
#define TMSG_ONTOP (TERMINAL_FIRST + 26)
#define INTERNET_ERROR_BASE 12000
#define ERR_FILE_EXISTS (INTERNET_ERROR_BASE + 224)
#define ERR_LOGON_FAILED (INTERNET_ERROR_BASE + 223)
#define ERR_NEWSGROUP_MISSING (INTERNET_ERROR_BASE + 411)
#define ERR_NO_ARTICLE (INTERNET_ERROR_BASE + 430)
#define ERR_NO_ARTICLE_NUMBER (INTERNET_ERROR_BASE + 423)
#define ERR_NO_ARTICLE_SELECTED (INTERNET_ERROR_BASE + 420)
#define ERR_NO_NEWSGROUP (INTERNET_ERROR_BASE + 412)
#define ERR_UNKNOWN_CODE_TYPE (INTERNET_ERROR_BASE + 225)
#define ERR_WSA_WAIT_TIMEOUT (INTERNET_ERROR_BASE + 258)
#define VOVER_BUILDNUMBER __VERSION__
#define __CAVOSTRMAXSTRING 256
#define __CAVOERRORSTRING "Cannot find string ("
#define RDT_FULL 1
#define RDT_TRANSFER 2
#define RDT_HIDDEN 8
#define SUCCESS 0
#define FAILURE -1
#define EDB 1000
#define EDB_SEEK (EDB + 1)
#define EDB_SKIP (EDB + 2)
#define EDB_GOTO (EDB + 3)
#define EDB_SETRELATION (EDB + 4)
#define EDB_USE (EDB + 5)
#define EDB_CREATEINDEX (EDB + 6)
#define EDB_SETORDER (EDB + 7)
#define EDB_SETINDEX (EDB + 8)
#define EDB_FIELDNAME (EDB + 9)
#define EDB_BADALIAS (EDB + 10)
#define EDB_DUPALIAS (EDB + 11)
#define EDB_SETFILTER (EDB + 12)
#define EDB_CYCLICREL (EDB + 13)
#define EDB_CREATETABLE (EDB + 14)
#define EDB_RDDNOTFOUND (EDB + 15)
#define EDB_FIELDINDEX (EDB + 17)
#define EDB_SELECT (EDB + 18)
#define EDB_SYMSELECT (EDB + 19)
#define EDB_TOTAL (EDB + 20)
#define EDB_RECNO (EDB + 21)
#define EDB_EXPRESSION (EDB + 22)
#define EDB_EXPR_WIDTH (EDB + 23)
#define EDB_DRIVERLOAD (EDB + 30)
#define EDB_PARAM (EDB + 31)
#define EDB_NOAREAS (EDB + 32)
#define EDB_NOMEM (EDB + 33)
#define EDB_NOFIELDS (EDB + 35)
#define EDB_BAD_ERROR_INFO (EDB + 36)
#define EDB_WRONGFIELDNAME (EDB + 37)
#define EDB_ORDDESTROY (EDB + 38)
#define EDB_NOINITFUNCTION (EDB + 39)
#define EDB_ERRORINIT (EDB + 40)
#define EDB_DBSTRUCT (EDB + 41)
#define EDB_NOTABLE (EDB + 50)
#define EDB_NOORDER (EDB + 51)
#define EDB_ASSERTION (EDB + 53)
#define DBI_ISDBF 1
#define DBI_CANPUTREC 2
#define DBI_GETHEADERSIZE 3
#define DBI_LASTUPDATE 4
#define DBI_GETDELIMITER 5
#define DBI_SETDELIMITER 6
#define DBI_GETRECSIZE 7
#define DBI_GETLOCKARRAY 8
#define DBI_TABLEEXT 9
#define DBI_READONLY 10
#define DBI_ISFLOCK 20
#define DBI_CHILDCOUNT 22
#define DBI_FILEHANDLE 23
#define DBI_FULLPATH 24
#define DBI_ISANSI 25
#define DBI_BOF 26
#define DBI_EOF 27
#define DBI_DBFILTER 28
#define DBI_FOUND 29
#define DBI_FCOUNT 30
#define DBI_LOCKCOUNT 31
#define DBI_VALIDBUFFER 32
#define DBI_ALIAS 33
#define DBI_GETSCOPE 34
#define DBI_LOCKOFFSET 35
#define DBI_SHARED 36
#define DBI_MEMOEXT 37
#define DBI_MEMOHANDLE 38

// duplicate define
#define DBI_BLOB_HANDLE 38
#define DBI_MEMOBLOCKSIZE 39
#define DBI_BLOB_INTEGRITY 40
#define DBI_CODEPAGE 41
#define DBI_BLOB_RECOVER 43
#define DBI_NEWINDEXLOCK 44
#define DBI_DB_VERSION 101
#define DBI_RDD_VERSION 102
#define DBI_RDD_LIST 103
#define DBI_MEMOFIELD 104
#define DBI_VO_MACRO_SYNTAX 105
#define DBI_USER 1000

#define DBOI_CONDITION 1
#define DBOI_EXPRESSION 2
#define DBOI_POSITION 3
#define DBOI_RECNO 4
#define DBOI_NAME 5
#define DBOI_NUMBER 6
#define DBOI_INDEXNAME 7
#define DBOI_INDEXEXT 8
// duplicate defines
#define DBOI_BAGNAME 7
#define DBOI_BAGEXT 8
#define DBOI_FULLPATH 20
#define DBOI_FILEHANDLE 21
#define DBOI_ISDESC 22
#define DBOI_ISCOND 23
#define DBOI_KEYTYPE 24
#define DBOI_KEYSIZE 25
#define DBOI_KEYCOUNT 26
#define DBOI_SETCODEBLOCK 27
#define DBOI_KEYDEC 28
#define DBOI_HPLOCKING 29
#define DBOI_LOCKOFFSET 35
#define DBOI_KEYADD 36
#define DBOI_KEYDELETE 37
#define DBOI_KEYVAL 38
#define DBOI_SCOPETOP 39
#define DBOI_SCOPEBOTTOM 40
#define DBOI_SCOPETOPCLEAR 41
#define DBOI_SCOPEBOTTOMCLEAR 42
#define DBOI_UNIQUE 43
#define DBOI_ORDERCOUNT 44
#define DBOI_CUSTOM 45
#define DBOI_SKIPUNIQUE 46
#define DBOI_KEYGOTO 47
#define DBOI_KEYSINCLUDED 48
#define DBOI_KEYNORAW 49
#define DBOI_OPTLEVEL 50
#define DBOI_KEYCOUNTRAW 51
#define DBOI_LOCK_ALL 100
#define DBOI_LOCK_FAIL 101
#define DBOI_HPLOCK_GATE 102
#define DBOI_USER 1000

#define TOPSCOPE 0
#define BOTTOMSCOPE 1

#define DBRI_DELETED 1
#define DBRI_LOCKED 2
#define DBRI_RECSIZE 3
#define DBRI_RECNO 4
#define DBRI_UPDATED 5
#define DBRI_BUFFPTR 6
#define DBRI_USER 1000

#define DBS_NAME 1
#define DBS_TYPE 2
#define DBS_LEN 3
#define DBS_DEC 4
#define DBS_ALIAS 5

#define DBS_BLOB_TYPE 102
#define DBS_BLOB_LEN 103
#define DBS_BLOB_POINTER 198
#define DBS_BLOB_DIRECT_TYPE 222
#define DBS_BLOB_DIRECT_LEN 223

#define DBS_STRUCT 998
#define DBS_PROPERTIES 999
#define DBS_USER 1000
#define BLOB_INFO_HANDLE 201
#define BLOB_FILE_RECOVER 202
#define BLOB_FILE_INTEGRITY 203
#define BLOB_OFFSET 204
#define BLOB_POINTER 205
#define BLOB_LEN 206
#define BLOB_TYPE 207
#define BLOB_EXPORT 208
#define BLOB_ROOT_UNLOCK 209
#define BLOB_ROOT_PUT 210
#define BLOB_ROOT_GET 211
#define BLOB_ROOT_LOCK 212
#define BLOB_IMPORT 213
#define BLOB_DIRECT_PUT 214
#define BLOB_DIRECT_GET 215
#define BLOB_GET 216
#define BLOB_DIRECT_EXPORT 217
#define BLOB_DIRECT_IMPORT 218
#define BLOB_NMODE 219
#define BLOB_EXPORT_APPEND 220
#define BLOB_EXPORT_OVERWRITE 221

#define BLOB_USER 1000
#define RDD_INFO                     100
#define _SET_MEMOBLOCKSIZE           101
#define _SET_DEFAULTRDD              102
#define _SET_MEMOEXT                 103
#define _SET_AUTOOPEN                104
#define _SET_AUTOORDER               105
#define _SET_HPLOCKING               106
#define _SET_NEWINDEXLOCK            107
#define _SET_AUTOSHARE               108
#define _SET_STRICTREAD              109
#define _SET_BLOB_CIRCULAR_ARRAY_REF 110
#define _SET_OPTIMIZE                111
#define _SET_FOXLOCK                 112
#define _SET_WINCODEPAGE             113
#define _SET_DOSCODEPAGE             114
#define RDD_INFO_MAX                 114
#define _SET_USER           (RDD_INFO + 100)
#define _SET_AXSLOADED      (_SET_USER + 1)

// defines used for the RL support in the DBFCDX driver
#define DBI_RL_AND          (DBI_USER + 1)
#define DBI_RL_CLEAR        (DBI_USER + 2)
#define DBI_RL_COUNT        (DBI_USER + 3)
#define DBI_RL_DESTROY      (DBI_USER + 4)
#define DBI_RL_EXFILTER     (DBI_USER + 5)
#define DBI_RL_GETFILTER    (DBI_USER + 6)
#define DBI_RL_HASMAYBE     (DBI_USER + 7)
#define DBI_RL_LEN          (DBI_USER + 8)
#define DBI_RL_MAYBEEVAL    (DBI_USER + 9)
#define DBI_RL_NEW          (DBI_USER + 10)
#define DBI_RL_NEWDUP       (DBI_USER + 11)
#define DBI_RL_NEWQUERY     (DBI_USER + 12)
#define DBI_RL_NEXTRECNO    (DBI_USER + 13)
#define DBI_RL_NOT          (DBI_USER + 14)
#define DBI_RL_OR           (DBI_USER + 15)
#define DBI_RL_PREVRECNO    (DBI_USER + 16)
#define DBI_RL_SET          (DBI_USER + 17)
#define DBI_RL_SETFILTER    (DBI_USER + 18)
#define DBI_RL_TEST         (DBI_USER + 19)



#define NEW_AREA 0
#define BUFF_SIZE 0x00008000
#define FO_CREATE 0x00001000
#ifndef MAXFILENAME
   #define MAXFILENAME 260
#endif
#define MAX_EXT_NAME 5
#define DB_MAXAREAS 1024
#define MAXDRIVERNAME 12
#define MAX_KEY_LEN 256
#define DBF_ANSI 0x04
#define DBF_VER 0x03
#define DBF_MEMO 0x80
#define DBF_DB4MEMO 0x88
#define DBF_PRODINDEX 0x01
#define DBF_MEMOS 0x02
#define DBF_ISDATABASE 0x04
#define DBF_OLE 0x80 
#define RDD_FUNCCOUNT (_SIZEOF(_RDDFUNCS)/4)
#define WAGNER_STRING (0)
#define WAGNER_OBJECT (2)
#define WAGNER_ARRAY (4)
#define WAGNER_FIXED (6)
#define WAGNER_FLOAT (8)
#define WAGNER_ARRAY_PAGE (10)
#define WAGNER_BINARY (0x40)
#define WAGNER_STATIC (0x80)
#define WAGNER_FORWARD (0xFFFD)
#define WAGNER_HAS_AXIT (0x80)
#define WAGNER_AXIT_CALLED (0x04)
#define WAGNER_OLDSPACE_STATE (0x02)
#define MAX_INST 10
#define F_ERROR PTR(_CAST,0xFFFFFFFF)
#define FERROR_FULL 256
#define FERROR_EOF 257
#define FERROR_PARAM 258
#define FS_SET 0
#define FS_RELATIVE 1
#define FS_END 2
#define FO_READ 0
#define FO_WRITE 1
#define FO_READWRITE 2
#define FO_COMPAT 0x00000000
#define FO_EXCLUSIVE 0x00000010
#define FO_DENYWRITE 0x00000020
#define FO_DENYREAD 0x00000030
#define FO_DENYNONE 0x00000040
#define FO_SHARED 0x00000040
#define FXO_WILD 0x00010000
#define FC_NORMAL 0x00000000
#define FC_READONLY 0x00000001
#define FC_HIDDEN 0x00000002
#define FC_SYSTEM 0x00000004
#define FC_ARCHIVED 0x00000020
#define FA_VOLUME 0x00000008
#define FA_DIRECTORY 0x00000010
#define FA_TEMPORARY 0x00000100
#define FA_COMPRESSED 0x00000800
#define FA_OFFLINE 0x00001000
#define F_NAME 1
#define F_SIZE 2
#define F_DATE 3
#define F_TIME 4
#define F_ATTR 5
#define F_LEN 5
#define PI 3.14159265358979323846
#define PI_2 1.57079632679489661923
#define PI_4 0.785398163397448309616
#define L2E 1.44269504088896340736
#define L2T 3.32192809488736234781
#define L10E 0.434294481903251827651
#define LG2 0.301029995663981195226
#define LN2 0.693147180559945309417
#define LN10 2.30258509299404568402
#define REAL4_EPSILON 1.192092896e-07
#define REAL4_MAX 3.402823466e+38
#define REAL8_EPSILON 2.2204460492503131e-016
#define REAL8_MAX 1.7976931348623158e+308
#define TICK_FREQUENCY 18.20647
#define ASC_BELL 7
#define ASC_BS 8
#define ASC_TAB 9
#define ASC_LF 10
#define ASC_FF 12
#define ASC_CR 13
#define ASC_SOFT_CR 141
#define ASC_EOF 26
#define ASC_ESC 27
#define ASC_BLANK 32
#define ASC_0 48
#define ASC_1 49
#define ASC_9 57
#define ASC_A 65
#define ASC_Z 90
//#define CRLF _CHR(ASC_CR) +_CHR(ASC_LF)
#define INI_GROUP_RUNTIME "CA-Visual Objects"
//#define NULL PTR(_CAST, 0L)
//#define NULL_PTR PTR(_CAST, 0L)
//#define NULL_ARRAY ARRAY(_CAST, 0L)
//#define NULL_OBJECT OBJECT(_CAST, 0L)
//#define NULL_DATE DATE(_CAST, 0L)
//#define NULL_CODEBLOCK CODEBLOCK(_CAST, 0L)
//#define NULL_STRING STRING(_CAST, 0L)
//#define NULL_PSZ PSZ(_CAST, 0L)
//#define NULL_SYMBOL SYMBOL(_CAST, 0)
#define KID_IN_AXIT 0x20000000
#define MAX_ALLOC 65527
#define _MAX_PATH 260
#define _MAX_DRIVE 3
#define _MAX_DIR 256
#define _MAX_FNAME 256
#define _MAX_EXT 256
#define MEMORY_COLLECT -1
#define MEMORY_SYSTEM_FREE 0
#define MEMORY_SYSTEM_MAX 1
#define MEMORY_DYNINFOFREE 2
#define MEMORY_DYNINFOMAX 3
#define MEMORY_KIDSTACK_SIZE 4
#define MEMORY_KIDSTACK_FREE 5
#define MEMORY_STACK_SIZE 6
#define MEMORY_STACK_FREE 7
#define MEMORY_MAXATOM 8
#define MEMORY_ACTIVATION 9
#define MEMORY_PUBLIC 10
#define MEMORY_PRIVAT 11
#define MEMORY_DYNINFOUSED 12
#define MEMORY_MEMTOTAL 13
#define MEMORY_DS_SIZE 14
#define MEMORY_CS_SIZE 15
#define MEMORY_REGISTEREXIT_COUNT 16
#define MEMORY_REGCOLLNOTIFYSTART_COUNT 17
#define MEMORY_REGCOLLNOTIFYEND_COUNT 18
#define MEMORY_REGISTERKID 19
#define MEMORY_REGISTERAXIT 20
#define MEMORY_COLLECTCOUNT 21
#define MEMORY_DYNINFOSIZE 22
#define MEMORY_RT_DGROUP 23
#define MEMORY_RT_DS 24
#define MEMORY_SS 25
#define MEMORY_DS 26
#define MEMORY_CS 27
#define MEMORY_SEQUENCE 28
#define MEMORY_STACKKID 29
#define MEMORY_SP 30
#define MEMORY_GLOBALSEL 31
#define MEMORY_FUNCTIONCOUNT 32
#define MEMORY_CLASSCOUNT 33
#define MEMORY_DB_DS 34
#define MEMORY_DB_DS_SIZE 35
#define MEMORY_WINDOWS_SYSTEMRESOURCES 100
#define MEMORY_WINDOWS_GDIRESOURCES 101
#define MEMORY_WINDOWS_USERRESOURCES 102
#define AMERICAN 1
#define ANSI 2
#define BRITISH 3
#define FRENCH 4
#define GERMAN 5
#define ITALIAN 6
#define JAPANESE 7
#define USA 8
#define JUL_BASE 1721060
#define CLASS_DEBUG_ALLOC 0x01
#define CLASS_DEBUG_INIT 0x02
#define CLASS_DEBUG_AXIT 0x04
#define CLASS_DEBUG_SEND 0x08
#define CLASS_DEBUG_IVARGET 0x10
#define CLASS_DEBUG_IVARPUT 0x20
#define CLASS_DEBUG_DECLARE 0x40
#define CLASS_DEBUG_UNDECL 0x80
#define CLASS_DEBUG_METHDECL 0x100
#define CLASS_DEBUG_NOIVARGET 0x200
#define CLASS_DEBUG_NOIVARPUT 0x400
#define CLASS_DEBUG_ALL 0xFFFFFFFF
#define _SET_EXACT 1
#define _SET_FIXED 2
#define _SET_DECIMALS 3
#define _SET_DATEFORMAT 4
#define _SET_EPOCH 5
#define _SET_PATH 6
#define _SET_DEFAULT 7
#define _SET_EXCLUSIVE 8
#define _SET_SOFTSEEK 9
#define _SET_UNIQUE 10
#define _SET_DELETED 11
#define _SET_CANCEL 12
#define _SET_DEBUG 13
#define _SET_TYPEAHEAD 14
#define _SET_COLOR 15
#define _SET_CURSOR 16
#define _SET_CONSOLE 17
#define _SET_ALTERNATE 18
#define _SET_ALTFILE 19
#define _SET_DEVICE 20
#define _SET_EXTRA 21
#define _SET_EXTRAFILE 22
#define _SET_PRINTER 23
#define _SET_PRINTFILE 24
#define _SET_MARGIN 25
#define _SET_BELL 26
#define _SET_CONFIRM 27
#define _SET_ESCAPE 28
#define _SET_INSERT 29
#define _SET_EXIT 30
#define _SET_INTENSITY 31
#define _SET_SCOREBOARD 32
#define _SET_DELIMITERS 33
#define _SET_DELIMCHARS 34
#define _SET_WRAP 35
#define _SET_MESSAGE 36
#define _SET_MCENTER 37
#define _SET_SCROLLBREAK 38
#define _SET_DIGITS 39
#define _SET_NETERR 40
#define _SET_HPLOCK 41
#define _SET_ANSI 44
#define _SET_YIELD 45
#define _SET_LOCKTRIES 46
#define _SET_DICT 98
#define _SET_INTL 99
#define _SET_COUNT 99
#define GC_TYPE_STACK 1
#define GC_TYPE_REGISTERKID 2
#define GC_ENTRY_MAX_STRSIZE 48
