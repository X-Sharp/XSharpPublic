#define IDM_EmptyShellMenu "EmptyShellMenu"
#define IDA_EmptyShellMenu "EmptyShellMenu"
#define IDM_EmptyShellMenu_File_ID 15001
#define IDM_EmptyShellMenu_File_Open_ID 15002
#define IDM_EmptyShellMenu_File_Print_Setup_ID 15004
#define IDM_EmptyShellMenu_File_Exit_ID 15006
#define IDM_EmptyShellMenu_Help_ID 15007
#define IDM_EmptyShellMenu_Help_Index_ID 15008
#define IDM_EmptyShellMenu_Help_Using_Help_ID 15009
#define IDM_EmptyShellMenu_Help_About_ID 15011
#define IDM_EmptyShellMenu_Help_dialogwindow1_ID 15012
#define IDM_StandardShellMenu "StandardShellMenu"
#define IDA_StandardShellMenu "StandardShellMenu"
#define IDM_StandardShellMenu_File_ID 15001
#define IDM_StandardShellMenu_File_Open_ID 15002
#define IDM_StandardShellMenu_File_Close_ID 15003
#define IDM_StandardShellMenu_File_Print_ID 15005
#define IDM_StandardShellMenu_File_Print_Setup_ID 15006
#define IDM_StandardShellMenu_File_Exit_ID 15008
#define IDM_StandardShellMenu_Edit_ID 15009
#define IDM_StandardShellMenu_Edit_Cut_ID 15010
#define IDM_StandardShellMenu_Edit_Copy_ID 15011
#define IDM_StandardShellMenu_Edit_Paste_ID 15012
#define IDM_StandardShellMenu_Edit_Insert_Record_ID 15014
#define IDM_StandardShellMenu_Edit_Delete_Record_ID 15015
#define IDM_StandardShellMenu_Edit_Go_To_Top_ID 15017
#define IDM_StandardShellMenu_Edit_Previous_ID 15018
#define IDM_StandardShellMenu_Edit_Next_ID 15019
#define IDM_StandardShellMenu_Edit_Go_To_Bottom_ID 15020
#define IDM_StandardShellMenu_View_ID 15021
#define IDM_StandardShellMenu_View_Form_ID 15022
#define IDM_StandardShellMenu_View_Table_ID 15023
#define IDM_StandardShellMenu_Window_ID 15024
#define IDM_StandardShellMenu_Window_Cascade_ID 15025
#define IDM_StandardShellMenu_Window_Tile_ID 15026
#define IDM_StandardShellMenu_Window_Close_All_ID 15027
#define IDM_StandardShellMenu_Help_ID 15028
#define IDM_StandardShellMenu_Help_Index_ID 15029
#define IDM_StandardShellMenu_Help_Context_Help_ID 15030
#define IDM_StandardShellMenu_Help_Using_Help_ID 15031
#define IDM_StandardShellMenu_Help_About_ID 15033
