﻿// $safeitemrootname$.vh
// Created by    : $username$
// Creation Date : $time$
// Created for   : $registeredorganization$
// WorkStation   : $machinename$


// Please note that XSharp supports both the Vulcan #define syntax as well as the Visual Objects define syntax:
// #define WM_USER 0x0400
// DEFINE WM_USER := 0x0400 AS DWORD