///////////////////////////////////////////////////////////////////////////
// VOOLEClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// OLE Classes library
//

#define BAS_NO 0
#define BAS_ONCE 1
#define BAS_ALWAYS 2
#define Unchecked 0
#define Checked 1
#define Gray 2
#define OFD_NAME 1
#define OFD_MEMBERID 2
#define OFD_INVOKE 3
#define OFD_PARAMS 4
#define OFD_OPTPARAMS 5
#define OFD_NAMEDARGS 6
#define OFD_PARAMDESC 7
#define OFD_RETDESC 8
#define OFD_LEN 8
#define TKIND_ENUM 0
#define TKIND_RECORD 1
#define TKIND_MODULE 2
#define TKIND_INTERFACE 3
#define TKIND_DISPATCH 4
#define TKIND_COCLASS 5
#define TKIND_ALIAS 6
#define TKIND_UNION 7
#define TKIND_MAX 8
#define VTS_I2 _CHR(0x02)
#define VTS_I4 _CHR(0x03)
#define VTS_R4 _CHR(0x04)
#define VTS_R8 _CHR(0x05)
#define VTS_CY _CHR(0x06)
#define VTS_DATE _CHR(0x07)
#define VTS_BSTRW _CHR(0x08)
#define VTS_DISPATCH _CHR(0x09)
#define VTS_SCODE _CHR(0x0A)
#define VTS_ERROR _CHR(0x0A)
#define VTS_BOOL _CHR(0x0B)
#define VTS_VARIANT _CHR(0x0C)
#define VTS_UNKNOWN _CHR(0x0D)
#define VTS_BSTRA _CHR(0x0E)
#define VTS_I1 _CHR(0x10)
#define VTS_UI1 _CHR(0x11)
#define VTS_UI2 _CHR(0x12)
#define VTS_UI4 _CHR(0x13)
#define VTS_I8 _CHR(0x14)
#define VTS_UI8 _CHR(0x15)
#define VTS_PI2 _CHR(0x42)
#define VTS_PI4 _CHR(0x43)
#define VTS_PR4 _CHR(0x44)
#define VTS_PR8 _CHR(0x45)
#define VTS_PCY _CHR(0x46)
#define VTS_PDATE _CHR(0x47)
#define VTS_PBSTR _CHR(0x48)
#define VTS_PDISPATCH _CHR(0x49)
#define VTS_PSCODE _CHR(0x4A)
#define VTS_PBOOL _CHR(0x4B)
#define VTS_PVARIANT _CHR(0x4C)
#define VTS_PUNKNOWN _CHR(0x4D)
#define VTS_PI1 _CHR(0x50)
#define VTS_PUI1 _CHR(0x51)
#define VTS_PUI2 _CHR(0x52)
#define VTS_PUI4 _CHR(0x53)
#define VTS_PI8 _CHR(0x54)
#define VTS_PUI8 _CHR(0x55)
#define VTS_AI2 _CHR(0x82)
#define VTS_AI4 _CHR(0x83)
#define VTS_AR4 _CHR(0x84)
#define VTS_AR8 _CHR(0x85)
#define VTS_ACY _CHR(0x86)
#define VTS_ADATE _CHR(0x87)
#define VTS_ABSTR _CHR(0x88)
#define VTS_ADISPATCH _CHR(0x89)
#define VTS_ASCODE _CHR(0x8A)
#define VTS_ABOOL _CHR(0x8B)
#define VTS_AVARIANT _CHR(0x8C)
#define VTS_AUNKNOWN _CHR(0x8D)
#define VTS_AI1 _CHR(0x90)
#define VTS_AUI1 _CHR(0x91)
#define VTS_AUI2 _CHR(0x92)
#define VTS_AUI4 _CHR(0x93)
#define VTS_AI8 _CHR(0x94)
#define VTS_AUI8 _CHR(0x95)
#define VT_VOBYREF 0x40
#define VT_VOARRAY 0x80
#define VT_VOMARKER 0xFF
