///////////////////////////////////////////////////////////////////////////
// VOSQLClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// SQL Classes library
//

#define _assert TRUE
#define __CAVO_SQL_TXN_READ_COMMITTED SQL_TXN_READ_COMMITTED
#define __CAVO_SQL_SIMULATE_CURSOR SQL_SC_TRY_UNIQUE
#define __CAVO_SQL_CURSOR_TYPE SQL_CURSOR_KEYSET_DRIVEN
#define __CAVO_SQL_CONCURRENCY SQL_CONCUR_ROWVER
#define __CAVO_SQL_ODBC_CURSORS SQL_CUR_USE_IF_NEEDED
#define __CAVO_SQL_MODE_READ_WRITE SQL_MODE_READ_WRITE
#define MAX_CONNECT_INFO_STRING 256
#define MAX_LONGVARCHAR 32000
#define MAX_LONGVARCHAR_EXT 100000
#define MAX_COLNAME_SIZE 40
#define SQL_RELOP_AND 1
#define SQL_RELOP_OR 2
#define SQL_RELOP_NOT 3
#define SQL_RELOP_OPENP 4
#define SQL_RELOP_CLOSEP 5
#define SQL_SC_UPD_AUTO 0
#define SQL_SC_UPD_CURSOR 1
#define SQL_SC_UPD_KEY 2
#define SQL_SC_UPD_VALUE 3
#define SQL_DATA_DELETE 1
#define SQL_DATA_BUFFER 2
#define SQL_DATA_NULL 3
#define SQL_LOGICAL_TRUE 0x31
#define SQL_LOGICAL_FALSE 0x30
#define SQL_BLANK_CHARACTER 0x20
#define __CAVOSTR_SQLCLASS__QE_LIC "IVC3.LIC"
#define __CAVOSTR_SQLCLASS__QE_PSWD "jys777JE04nN13Ef52eR4x3b"
#define __CAVOSTR_SQLCLASS__IS_NULL " IS NULL"
#define __CAVOSTR_SQLCLASS__NULL " NULL"
#define __CAVOSTR_SQLCLASS__1_QUOTE "'"
#define __CAVOSTR_SQLCLASS__2_QUOTE "''"
#define __CAVOSTR_SQLCLASS__SELECT "select "
#define __CAVOSTR_SQLCLASS__FROM " from "
#define __CAVOSTR_SQLCLASS__UPDATE "update "
#define __CAVOSTR_SQLCLASS__SET " set "
#define __CAVOSTR_SQLCLASS__CURR_OF " where current of "
#define __CAVOSTR_SQLCLASS__WHERE " where "
#define __CAVOSTR_SQLCLASS__AND " and "
#define __CAVOSTR_SQLCLASS__DEL_FROM "delete from "
#define __CAVOSTR_SQLCLASS__INS_INTO "insert into "
#define __CAVOSTR_SQLCLASS__VALUES ") values ("
#define __CAVOSTR_SQLCLASS__ORDER_BY " order by "
#define __CAVOSTR_SQLCLASS__DSN "DSN="
#define __CAVOSTR_SQLCLASS__UID "UID="
#define __CAVOSTR_SQLCLASS__PWD "PWD="
#define __CAVOSTR_SQLCLASS__EQ_NULL " = NULL"
#define __CAVOSTR_SQLCLASS__EQ " ="
#define SQL_TYPE_UNKNOWN -9999
