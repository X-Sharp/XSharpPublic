///////////////////////////////////////////////////////////////////////////
// VOGUIClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// GUI Classes library
//

#define __WCCustomControlClass "_VOCustomControl"
#define GBSSBLEFT 1
#define GBSSBMIDDLE 2
#define GBSSBRIGHT 3
#define ssBlockSelection 3
#define ssExtendedSelection 2
#define ssNoSelection 0
#define ssSingleSelection 1
#define __WCGBNotifyWindowClass "GBNotifyContext"
#define __WCDocAppWindowClass "DocAppWindow"
#define WM_DRAGSELECT 0x022E
#define WM_QUERYDROPOBJECT 0x022B
#define FSEL_ALL 0
#define FSEL_END 3
#define FSEL_HOME 2
#define FSEL_TRIM 1
#define FSEL_TRIMEND 4
#define MAX_FMTSTRING_LEN 4096
#define OVERWRITE_ALWAYS 2
#define OVERWRITE_NEVER 0
#define OVERWRITE_ONKEY 1
#define SCRMODE_FULL 0
#define SCRMODE_NO 2
#define SCRMODE_PART 1
#define DEFAULT_STRING_TEMPL_SIZE 128
#define INSIDEFORMBORDER 5
#define MIN_DATAWINDOWWIDTH 50
#define HDCANTOPENFILE 1
#define HDINVALIDKEY 3
#define HDOK 0
#define HDOUTOFMEMORY 2
#define HDUNKNOWN 4
#define Max_Wait 2000
#define __WCMMContWindowClass "_VOMMContainer"
#define MM_AVI 2
#define MM_BMP 1
#define MM_UNKNOWN 0
#define MM_WAV 3
#define OLEPROP_ACTIVATEONDBLCLK 0x00000002L
#define OLEPROP_ALLOWDOCVIEW 0x00000040L
#define OLEPROP_ALLOWINPLACE 0X00000001L
#define OLEPROP_ALLOWRESIZE 0x00000004L
#define OLEPROP_AUTOSIZEONCREATE 0x00000008L
#define OLEPROP_ISACTIVE 0x00000020L
#define OLEPROP_READONLY 0x00000010L
#define USERclassTYPE_APPNAME 3
#define USERclassTYPE_FULL 1
#define USERclassTYPE_SHORT 2
#define DROPEFFECT_COPY 1
#define DROPEFFECT_LINK 4
#define DROPEFFECT_MOVE 2
#define DROPEFFECT_NONE 0
#define IDM_OLE_CONVERT 57343
#define IDM_OLE_VERB_FIRST 57280
#define IDM_OLE_VERB_LAST 57342
#define MAX_NAME 260
#define OLE_DDEVENT_DRAGENTER 1
#define OLE_DDEVENT_DRAGLEAVE 2
#define OLE_DDEVENT_DRAGOVER 3
#define OLE_DDEVENT_DROP 4
#define OLECMDEXECOPT_DODEFAULT 0
#define OLECMDEXECOPT_DONTPROMPTUSER 2,
#define OLECMDEXECOPT_PROMPTUSER 1
#define OLECMDEXECOPT_SHOWHELP 3
#define OLECMDID_CLEARSELECTION 18
#define OLECMDID_COPY 12
#define OLECMDID_CUT 11
#define OLECMDID_GETZOOMRANGE 20
#define OLECMDID_HIDETOOLBARS 24
#define OLECMDID_NEW 2
#define OLECMDID_OPEN 1
#define OLECMDID_PAGESETUP 8
#define OLECMDID_PASTE 13
#define OLECMDID_PASTESPECIAL 14
#define OLECMDID_PRINT 6
#define OLECMDID_PRINTPREVIEW 7
#define OLECMDID_PROPERTIES 10
#define OLECMDID_REDO 16
#define OLECMDID_REFRESH 22
#define OLECMDID_SAVE 3
#define OLECMDID_SAVEAS 4
#define OLECMDID_SAVECOPYAS 5
#define OLECMDID_SELECTALL 17
#define OLECMDID_SETDOWNLOADSTATE 29
#define OLECMDID_SETPROGRESSMAX 25
#define OLECMDID_SETPROGRESSPOS 26
#define OLECMDID_SETPROGRESSTEXT 27
#define OLECMDID_SETTITLE 28
#define OLECMDID_SPELL 9
#define OLECMDID_STOP 23
#define OLECMDID_STOPDOWNLOAD 30
#define OLECMDID_UNDO 15
#define OLECMDID_UPDATECOMMANDS 21
#define OLECMDID_ZOOM 19
#define CAPABILITY_NOT_AVAILABLE 0xFFFFFFFF
#define CCHBINNAME 24
#define CCHPAPERNAME 64
#define EM_SETTYPOGRAPHYOPTIONS (WM_USER + 202)
#define RICHTAB_CENTER 0x01000000
#define RICHTAB_DECIMAL 0x03000000
#define RICHTAB_NORMAL 0x00000000
#define RICHTAB_RIGHT 0x02000000
#define RICHTAB_WORDBAR 0x04000000
#define TO_ADVANCEDTYPOGRAPHY 1
#define TO_SIMPLELINEBREAK 2
#define RICHEDIT_CLASS "RichEdit20A"
#define TBL_CHILD 0
#define TBL_SHELL 1
#define TBL_SHELLBAND 2
#define __WCShellWindowClass "ShellWindow"
#define BFFM_ENABLEOK (WM_USER + 101)
#define BFFM_INITIALIZED 1
#define BFFM_SELCHANGED 2
#define BFFM_SETSELECTION (WM_USER + 102)
#define BFFM_SETSTATUSTEXT (WM_USER + 100)
#define BIF_BROWSEFORCOMPUTER 0x1000
#define BIF_BROWSEFORPRINTER 0x2000
#define BIF_BROWSEINCLUDEFILES 0x4000
#define BIF_DONTGOBELOWDOMAIN 0x0002
#define BIF_RETURNFSANCESTORS 0x0008
#define BIF_RETURNONLYFSDIRS 0x0001
#define BIF_STATUSTEXT 0x0004
#define SB_SETICON (WM_USER+15)
#define SBT_TOOLTIPS 0x0800
#define iPageBorder 2
#define ECM_FIRST 0x1500
#define EM_SETCUEBANNER (ECM_FIRST + 1)
#define EM_GETCUEBANNER (ECM_FIRST + 2)
#define EM_SHOWBALLOONTIP (ECM_FIRST + 3)
#define EM_HIDEBALLOONTIP (ECM_FIRST + 4)
#define TTI_NONE 0
#define TTI_INFO 1
#define TTI_WARNING 2
#define TTI_ERROR 3
#define I_IMAGENONE (-2)
#define RB_MAXIMIZEBAND (WM_USER + 31)
//#define TB_GETMAXSIZE WM_USER + 83
#define __WCTopAppWindowClass "TopAppWindow"
#define API_WINDOW_HDC 2
#define API_WINDOW_HWND 0
#define btNoBorder 0
#define btNonSizingBorder 2
#define btSizingBorder 1
#define Color_EndColors COLOR_BTNHIGHLIGHT
#define CONTAINER_CLASS "Ca_Container32"
#define FONTFAMILY_ANY 1000
#define FONTFAMILY_DECORAT 1005
#define FONTFAMILY_MODERN 1003
#define FONTFAMILY_ROMAN 1001
#define FONTFAMILY_SCRIPT 1004
#define FONTFAMILY_SWISS 1002
#define gbaAlignCenter 2
#define gbaAlignLeft 0
#define gbaAlignRight 1
#define gblButton 3
#define gblCaption 0
#define gblColButton 4
#define gblColCaption 2
#define gblHiText 5
#define gblText 1
#define GBNFY_CLOSE 13
#define GBNFY_COMPLETION 7
#define GBNFY_DEFERNOTIFY 11
#define GBNFY_DODELETE 6
#define GBNFY_DOGOEND 4
#define GBNFY_DOGOTOP 3
#define GBNFY_DONEWROW 5
#define GBNFY_DOSKIP 2
#define GBNFY_FIELDCHANGE 8
#define GBNFY_FILECHANGE 9
#define GBNFY_INTENTTOMOVE 10
#define GBNFY_PROCESSNOTIFY 12
#define GBNFY_RECORDCHANGE 1
#define GBNFY_VIEWASBROWSER 15
#define GBNFY_VIEWASFORM 16
#define GBNFY_VIEWSWITCH 14
#define gbsControl2d 2
#define gbsControl3d 1
#define gbsEdit 3
#define gbsReadOnly 0
#define LBAddString 1L
#define LBInsertString 2L
#define LBDeleteString 3L
#define LBFindString 4L
#define LBGetCount 5L
#define LBGetCurSel 6L
#define LBGetText 7L
#define LBGetTextLen 8L
#define LBResetContent 9L
#define LBSetCurSel 10L
#define LBFindStringExact 11L
#define MAX_LEN 4096
#define OFN_BIDIDIALOG 0X80000000
#define PICTYPE_CHAR 3
#define PICTYPE_DATE 2
#define PICTYPE_LOGICAL 5
#define PICTYPE_MEMO 4
#define PICTYPE_NUMERIC 1
#define PICTYPE_UNKNOWN 0
#define WCCartesianCoordinates TRUE
#define WCWindowsCoordinates FALSE
#define ID_FIRSTWCHELPID 0xFFFD
#define ID_WCHELP 0xFFFF
#define ID_WCHELPOFF 0xFFFD
#define ID_WCHELPON 0xFFFE
#define IDT_3DAREACHART 56
#define IDT_3DBARCHART 57
#define IDT_3DCOLUMNAREACHART 59
#define IDT_3DCOLUMNCHART 58
#define IDT_3DFRAME 86
#define IDT_3DLINECHART 60
#define IDT_3DPIECHART 61
#define IDT_3DSURFACECHART 62
#define IDT_ADDTEXT 25
#define IDT_ARC 73
#define IDT_AREACHART 49
#define IDT_ARROW 69
#define IDT_BACK 84
#define IDT_BARCHART 50
#define IDT_BOLD 08
#define IDT_BORDERLOW 29
#define IDT_BORDERRECT 28
#define IDT_BULLETLIST 104
#define IDT_BUTTON 45
#define IDT_CALC 89
#define IDT_CALCULATE 48
#define IDT_CENTER 22
#define IDT_CENTERTAB 116
#define IDT_CENTERTEXT 26
#define IDT_CHARTFORMAT 66
#define IDT_CLOSE 03
#define IDT_COLOR 85
#define IDT_COLUMNCHART 51
#define IDT_COLUMNFORMAT 107
#define IDT_COLUMNLINECHART 64
#define IDT_COLUMNSTOCKCHART 65
#define IDT_COMMA 18
#define IDT_COPY 31
#define IDT_CROSSOUT 11
#define IDT_CURRENCY 16
#define IDT_CUSTOMBITMAP 132
#define IDT_CUT 101
#define IDT_DECIMALMINUS 20
#define IDT_DECIMALPLUS 19
#define IDT_DECIMALTAB 118
#define IDT_DELETE 121
#define IDT_DISKETTEIO 125
#define IDT_EDITCHART 67
#define IDT_EDITPOINT 80
#define IDT_ELLIPSE 72
#define IDT_ENDREC 130
#define IDT_ENVELOPE 111
#define IDT_FILLEDARC 77
#define IDT_FILLEDELLIPSE 76
#define IDT_FILLEDPOLYGON 78
#define IDT_FILLEDRECTANGLE 75
#define IDT_FIND 126
#define IDT_FRAME 108
#define IDT_FREEHAND 70
#define IDT_FRONT 83
#define IDT_FUNCTION 88
#define IDT_GOMACRO 90
#define IDT_GRAPH 110
#define IDT_GROUP 81
#define IDT_HELP 120
#define IDT_INDENT 106
#define IDT_ITALIC 09
#define IDT_JUSTIFY 24
#define IDT_LEFT 21
#define IDT_LEFTTAB 115
#define IDT_LIGHTSHADING 30
#define IDT_LINE 68
#define IDT_LINECHART 53
#define IDT_LOCK 40
#define IDT_MAIL 123
#define IDT_NEW 100
#define IDT_NEWMACRO 87
#define IDT_NEWSHEET 01
#define IDT_NEXTREC 128
#define IDT_NUMBERLIST 103
#define IDT_OBJECT 109
#define IDT_OPEN 02
#define IDT_OUTLINESYMBOL 41
#define IDT_PAGEFIT 114
#define IDT_PAGELAYOUT 112
#define IDT_PAGENORMAL 113
#define IDT_PARAGRAPH 119
#define IDT_PASTE 102
#define IDT_PASTEFORMAT 32
#define IDT_PASTEVALUE 33
#define IDT_PAUSEMACRO 99
#define IDT_PERCENT 17
#define IDT_PICTURE 46
#define IDT_PIECHART 54
#define IDT_POLYGON 74
#define IDT_PREVIEW 06
#define IDT_PREVREC 127
#define IDT_PRINT 05
#define IDT_RADARCHART 63
#define IDT_RECORDMACRO 97
#define IDT_RECTANGLE 71
#define IDT_REPEAT 35
#define IDT_RESETMACRO 96
#define IDT_RIGHT 23
#define IDT_RIGHTTAB 117
#define IDT_RUNMACRO 94
#define IDT_SAVE 04
#define IDT_SCATTERCHART 55
#define IDT_SCROLLMINUS 43
#define IDT_SCROLLPLUS 44
#define IDT_SELECTCELL 42
#define IDT_SELECTOBJECT 79
#define IDT_SEPARATOR 00
#define IDT_SIZEMINUS 13
#define IDT_SIZEPLUS 12
#define IDT_SKIPMACRO 95
#define IDT_SORTATOZ 38
#define IDT_SORTZTOA 39
#define IDT_SPELLCHECK 47
#define IDT_STACKCHART 52
#define IDT_STARTREC 129
#define IDT_STEPMACRO 91
#define IDT_STOPMACRO 98
#define IDT_SUBSCRIPT 15
#define IDT_SUM 07
#define IDT_SUPERSCRIPT 14
#define IDT_TABLE 27
#define IDT_TIME 122
#define IDT_TRACEINMACRO 93
#define IDT_TRACEOUTMACRO 92
#define IDT_TUTORIAL 124
#define IDT_UNDERLINE 10
#define IDT_UNDO 34
#define IDT_UNGROUP 82
#define IDT_UNINDENT 105
#define IDT_VFORM 132
#define IDT_VGBROWSE 131
#define IDT_ZOOMIN 36
#define IDT_ZOOMOUT 37
#define __WCWndAppWindowClass "WndAppWindow"
#define ARRANGEASICONS 0
#define ARRANGECASCADE 1
#define ARRANGETILE 2
#define ARRANGETILEHORIZONTAL 3
#define ARRANGETILEVERTICAL ARRANGETILE
#define BITMAPFORMAT 1
#define BLOCKDECREMENT 5
#define BLOCKINCREMENT 1
#define BMP_2DTRANSPARENT LR_LOADTRANSPARENT
#define BMP_3DTRANSPARENT LR_LOADMAP3DCOLORS
#define BMP_OPAQUE 0
#define BOXABORTRETRYIGNORE 2
#define BOXDROPDOWN 1
#define BOXDROPDOWNLIST 2
#define BOXICONASTERISK 0x40
#define BOXICONEXCLAMATION 0x30
#define BOXICONHAND 0x10
#define BOXICONQUESTIONMARK 0X20
#define BOXREPLYABORT 0
#define BOXREPLYCANCEL 1
#define BOXREPLYIGNORE 2
#define BOXREPLYNO 3
#define BOXREPLYOKAY 4
#define BOXREPLYRETRY 5
#define BOXREPLYYES 6
#define BOXREPLYCLOSE    7
#define BOXREPLYTRYAGAIN 8
#define BOXREPLYCONTINUE 9

#define BOXRTLREADING 0x0400
#define BOXSIMPLE 0
#define BOXSORTEDASCENDING 0
#define BOXSORTEDDESCENDING 1
#define BOXUNSORTED 2
#define BRUSHBLACK 7
#define BRUSHCLEAR 6
#define BRUSHDARK 1
#define BRUSHHOLLOW 5
#define BRUSHLIGHT 3
#define BRUSHMEDIUM 2
#define BRUSHWHITE 4
#define BUTTONCONTROL 8
#define BUTTONLEFT 1
#define BUTTONMIDDLE 16
#define BUTTONOKAY 0
#define BUTTONOKAYCANCEL 1
#define BUTTONRETRYCANCEL 5
#define BUTTONRIGHT 2
#define BUTTONSHIFT 4
#define BUTTONYESNO 4
#define BUTTONYESNOCANCEL 3
#define ButtonX1 0x0020
#define ButtonX2 0x0040
#define XBUTTON1 0x0001
#define XBUTTON2 0x0002
#define COLORBLACK 0
#define COLORBLUE 1
#define COLORCYAN 3
#define COLORGREEN 2
#define COLORMAGENTA 5
#define COLORRED 4
#define COLORWHITE 7
#define COLORYELLOW 6
#define EDITAUTOHSCROLL 0x00000080L
#define EDITAUTOVSCROLL 0x00000040L
#define EDITBORDERED 0x00800000L
#define EDITCENTER 0x00000001L
#define EDITHSCROLL 0x00100000L
#define EDITLEFT 0x00000000L
#define EDITLOWERCASE 0x00000010L
#define EDITMULTILINE 0x00000004L
#define EDITNOHIDESEL 0x00000100L
#define EDITOEMCONVERT 0x00000400L
#define EDITPASSWORD 0x00000020L
#define EDITREADONLY 0x00000800L
#define EDITRIGHT 0x00000002L
#define EDITUPPERCASE 0x00000008L
#define EDITVSCROLL 0x00200000L
#define EDITWANTRETURN 0x00001000L
#define EXECNORMAL 0
#define EXECWHILEEVENT 1
#define FONTANY 1
#define FONTDECORATIVE 0
#define FONTMODERN 2
#define FONTMODERN10 1
#define FONTMODERN12 2
#define FONTMODERN8 0
#define FONTROMAN 3
#define FONTROMAN10 4
#define FONTROMAN12 5
#define FONTROMAN14 6
#define FONTROMAN18 7
#define FONTROMAN24 8
#define FONTROMAN8 3
#define FONTSCRIPT 4
#define FONTSWISS 5
#define FONTSWISS10 10
#define FONTSWISS12 11
#define FONTSWISS14 12
#define FONTSWISS18 13
#define FONTSWISS24 14
#define FONTSWISS8 9
#define FONTSYSTEM8 15
#define FORMATBITMAP 1
#define FORMATTEXT 0
#define FT_CENTERED 1
#define FT_LEFTALIGN 0
#define FT_RIGHTALIGN 2
#define HATCHDIAGONAL135 3
#define HATCHDIAGONAL45 1
#define HATCHDIAGONALCROSS 6
#define HATCHHORIZONTAL 4
#define HATCHORTHOGONALCROSS 5
#define HATCHSOLID 0
#define HATCHVERTICAL 2
#define HELPCONTROL 1
#define HELPMENU 0
#define HELPWINDOW 2
#define HELPINFO 3
#define HM_GENERAL 1
#define HM_MOUSE 2
#define HM_NONE 3
#define ICONASTERISK 4
#define ICONEXCLAMATION 3
#define ICONHAND 1
#define ICONQUESTIONMARK 2
#define ICONSTANDARD 5
#define IDLEEXEC FALSE
#define IDLEINIT TRUE
#define IPCITEMNOTFOUND 3
#define IPCOUTOFMEMORY 1
#define IPCSERVERNOTFOUND 0
#define IPCTOPICNOTFOUND 2
#define KEYALT 0X12
#define KEYARROWDOWN 0X28
#define KEYARROWLEFT 0X25
#define KEYARROWRIGHT 0X27
#define KEYARROWUP 0X26
#define KEYBACKSPACE 0X08
#define KEYCANCEL 0X03
#define KEYCAPSLOCK 0X14
#define KEYCONTROL 0X11
#define KEYDELETE 0X2E
#define KEYEND 0X23
#define KEYENTER 0X0D
#define KEYESCAPE 0X1B
#define KEYF1 0X70
#define KEYF10 0X79
#define KEYF11 0X7A
#define KEYF12 0X7B
#define KEYF13 0X7C
#define KEYF14 0X7D
#define KEYF15 0X7E
#define KEYF16 0X7F
#define KEYF2 0X71
#define KEYF3 0X72
#define KEYF4 0X73
#define KEYF5 0X74
#define KEYF6 0X75
#define KEYF7 0X76
#define KEYF8 0X77
#define KEYF9 0X78
#define KEYHOME 0X24
#define KEYINSERT 0X2D
#define KEYNUMLOCK 0X90
#define KEYPAGEDOWN 0X22
#define KEYPAGEUP 0X21
#define KEYPAUSE 0X13
#define KEYPRINT 0X2A
#define KEYRETURN 0X0D
#define KEYSHIFT 0X10
#define KEYSPACE 0X20
#define KEYTAB 0X09
#define LBOXDISABLENOSCROLL 0x1000L
#define LBOXEXTENDEDSEL 0x0800L
#define LBOXHASSTRINGS 0x0040L
#define LBOXMULTICOLUMN 0x0200L
#define LBOXMULTIPLESEL 0x0008L
#define LBOXNOINTEGRALHEIGHT 0x0100L
#define LBOXNOREDRAW 0x0004L
#define LBOXNOTIFY 0x0001L
#define LBOXOWNERDRAWFIXED 0x0010L
#define LBOXOWNERDRAWVARIABLE 0x0020L
#define LBOXSORT 0x0002L
#define LBOXUSETABSTOPS 0x0080L
#define LBOXWANTKEYBOARDINPUT 0x0400L
#define LINECLEAR 5
#define LINEDASHDOT 3
#define LINEDASHDOTDOT 4
#define LINEDASHED 1
#define LINEDOTTED 2
#define LINESOLID 0
#define LV_GNIABOVE LVNI_ABOVE
#define LV_GNIBELOW LVNI_BELOW
#define LV_GNIBYITEM LVNI_ALL
#define LV_GNILEFT LVNI_TOLEFT
#define LV_GNIRIGHT LVNI_TORIGHT
#define LV_SEEKDOWN 2
#define LV_SEEKTEXT 0
#define LV_SEEKUP 3
#define LV_SEEKVALUE 1
#define MENUSEPARATOR -1
#define MESSAGECONTROL 3
#define MESSAGEERROR 4
#define MESSAGEMENU 2
#define MESSAGEPERMANENT 1
#define MESSAGEPRIORITY 3
#define MESSAGETRANSIENT 2
//#define OFF FALSE
//#define ON TRUE
#define PAINTFILL 0
#define PAINTFRAME 2
#define PAINTINVERT 1
#define PITCHFIXED 1
#define PITCHVARIABLE 2
#define PM_ALIGNCENTER TPM_CENTERALIGN
#define PM_ALIGNLEFT TPM_LEFTALIGN
#define PM_ALIGNRIGHT TPM_RIGHTALIGN
#define PM_LEFTBUTTON TPM_LEFTBUTTON
#define PM_RIGHTBUTTON TPM_RIGHTBUTTON
#define POINTERAPPSTARTING 7
#define POINTERARROW 6
#define POINTERCROSSHAIRS 0
#define POINTERFOURARROW 3
#define POINTERHOURGLASS 5
#define POINTERIBEAM 1
#define POINTERICON 2
#define POINTERUPARROW 4
#define PRINTERERRORFATALDEVICEERROR 0
#define PRINTERERRORGENERALERROR 4
#define PRINTERERRORNODISKSPACE 2
#define PRINTERERRORNOMEMSPACE 3
#define PRINTERERRORUSERABORT 1
#define REGIONBORDER 6
#define REGIONCANVAS 0
#define REGIONCAPTION 1
#define REGIONCLOSE 9
#define REGIONMAXBOX 4
#define REGIONMENUBAR 8
#define REGIONMINBOX 3
#define REGIONSIZEBOX 2
#define REGIONSYSTEMMENUBOX 5
#define REGIONUNKNOWN 7
#define REGWB_ISDELIMITER WB_ISDELIMITER
#define REGWB_LEFT WB_LEFT
#define REGWB_LEFTBREAK WB_LEFTBREAK
#define REGWB_MOVEWORDLEFT WB_MOVEWORDLEFT
#define REGWB_MOVEWORDRIGHT WB_MOVEWORDRIGHT
#define REGWB_RIGHT WB_RIGHT
#define REGWB_RIGHTBREAK WB_RIGHTBREAK
#define REOPT_AUTOHSCROLL ECO_AUTOHSCROLL
#define REOPT_AUTOVSCROLL ECO_AUTOVSCROLL
#define REOPT_AUTOWORD ECO_AUTOWORDSELECTION
#define REOPT_NOHIDESEL ECO_NOHIDESEL
#define REOPT_READONLY ECO_READONLY
#define REOPT_SAVESEL ECO_SAVESEL
#define REOPT_SELBAR ECO_SELECTIONBAR
#define REOPT_VERTICAL ECO_VERTICAL
#define REOPT_WANTRETURN ECO_WANTRETURN
#define REPARA_BULLET PFN_BULLET
#define REPARA_CENTER PFA_CENTER
#define REPARA_LEFT PFA_LEFT
#define REPARA_NUMBER 0
#define REPARA_RIGHT PFA_RIGHT
#define RESEL_EMPTY SEL_EMPTY
#define RESEL_MULTICHAR SEL_MULTICHAR
#define RESEL_MULTIOBJECT SEL_MULTIOBJECT
#define RESEL_OBJECT SEL_OBJECT
#define RESEL_TEXT SEL_TEXT
#define RESTR_RTF SF_RTF
#define RESTR_TEXT SF_TEXT
#define ROPBACKGROUND 1
#define ROPINVERT 2
#define ROPOVERWRITE 0
#define ROPXOR 3
#define SBITEMFLAT SBT_NOBORDERS
#define SBITEMRAISED SBT_POPOUT
#define SBITEMSUNKEN 0
#define SC_MASK 0xFFF0
#define SCROLLEND 0
#define SCROLLHORIZONTAL 4
#define SCROLLTHUMBDRAG 3
#define SCROLLTOBOTTOMRIGHT 7
#define SCROLLTOTOPLEFT 6
#define SCROLLVERTICAL 5
#define SHOWCENTERED 3
#define SHOWICONIZED 2
#define SHOWINACTIVE 4
#define SHOWNORMAL 0
#define SHOWZOOMED 1
#define SPLIT_COLORBAR SPLTCOLOR_BAR
#define SPLIT_COLORFRAME SPLTCOLOR_BARFRAME
#define SPLIT_COLORWINDOW SPLTCOLOR_WINDOW
#define SPLIT_HORZALIGN SWS_HALIGN
#define SPLIT_VERTALIGN SWS_VALIGN
#define STATUSCAPSLOCK 2
#define STATUSINSERT 0
#define STATUSKEYBOARD 4
#define STATUSMEMORY 3
#define STATUSMESSAGE 5
#define STATUSNUMLOCK 3
#define STATUSPAIR 2
#define STATUSSCROLLLOCK 1
#define STATUSTIME 1
#define STRINGFORMAT 0
#define SYSMENU_Mask 0xF000
//#define TB_BOTTOM 1
#define TB_CONCAVE 1
#define TB_CONVEX 2
#define TB_DEFSTRING "toolbar_defstring"
#define TB_DISABLE 0
#define TB_ENABLE 3
#define TB_FLOATING 4
#define TB_ICONONLY 1
//#define TB_LEFT 2
#define TB_NORMAL 1
#define TB_NOSTRING "toolbar_nostring"
#define TB_PLAIN 0
#define TB_RIGHT 3
#define TB_SELECT 2
#define TB_TEXTANDICON 2
#define TB_TEXTONLY 0
//#define TB_TOP 0
#define TEXTCENTERED 2
#define TEXTLEFTALIGN 0
#define TEXTRIGHTALIGN 1
#define TWIPSCONVERSION 20
#define UNITDECREMENT 4
#define UNITINCREMENT 2
#define WC_ctrl_mask 0XE000
#define WEIGHTHEAVY 2
#define WEIGHTLIGHT 1
#define WEIGHTNORMAL 0
#define WINDOWNOBORDER 0
#define WINDOWNONSIZINGBORDER 2
#define WINDOWSIZINGBORDER 1
#define WM_WCHelp 0XBFFF
#define TRAYTIP_LENGTH_SHELLORIGINAL 64
#define TRAYTIP_LENGTH_SHELL5 128
#define OA_LEFT 1
#define OA_LEFT_AUTOSIZE 5
#define OA_NO 0
#define OA_RIGHT 3
#define OA_RIGHT_AUTOSIZE 7
#define OA_TOP 2
#define OA_TOP_AUTOSIZE 6
#define OA_BOTTOM 4
#define OA_BOTTOM_AUTOSIZE 8
#define OA_CENTER 9
#define OA_FULL_SIZE 10
#define OA_HEIGHT 0b0000000110000000
#define OA_PHEIGHT 0b0000001110000000
#define OA_WIDTH 0b0000010010000000
#define OA_PWIDTH 0b0000110010000000
#define OA_WIDTH_HEIGHT (OA_WIDTH | OA_HEIGHT)
#define OA_WIDTH_PHEIGHT (OA_WIDTH | OA_PHEIGHT)
#define OA_PWIDTH_HEIGHT (OA_PWIDTH | OA_HEIGHT)
#define OA_PWIDTH_PHEIGHT (OA_PWIDTH | OA_PHEIGHT)
#define OA_HEIGHT_WIDTH OA_WIDTH_HEIGHT
#define OA_HEIGHT_PWIDTH OA_PWIDTH_HEIGHT
#define OA_PHEIGHT_WIDTH OA_WIDTH_PHEIGHT
#define OA_PHEIGHT_PWIDTH OA_PWIDTH_PHEIGHT
#define OA_X 0b0100000010000000
#define OA_Y 0b0001000010000000
#define OA_PX 0b1100000010000000
#define OA_PY 0b0011000010000000
#define OA_PX_HEIGHT (OA_PX | OA_HEIGHT)
#define OA_PX_PHEIGHT (OA_PX | OA_PHEIGHT)
#define OA_PX_WIDTH (OA_PX | OA_WIDTH)
#define OA_PX_PWIDTH (OA_PX | OA_PWIDTH)
#define OA_PX_PWIDTH_HEIGHT (OA_PX | OA_PWIDTH | OA_HEIGHT)
#define OA_PX_WIDTH_HEIGHT (OA_PX | OA_WIDTH | OA_HEIGHT)
#define OA_PX_PWIDTH_PHEIGHT (OA_PX | OA_PWIDTH | OA_PHEIGHT)
#define OA_PY_HEIGHT (OA_PY | OA_HEIGHT)
#define OA_PY_PHEIGHT (OA_PY | OA_PHEIGHT)
#define OA_PY_WIDTH (OA_PY | OA_WIDTH)
#define OA_PY_PWIDTH (OA_PY | OA_PWIDTH)
#define OA_PY_WIDTH_HEIGHT (OA_PY | OA_WIDTH | OA_HEIGHT)
#define OA_PY_WIDTH_PHEIGHT (OA_PY | OA_WIDTH | OA_PHEIGHT)
#define OA_PY_PWIDTH_HEIGHT (OA_PY | OA_PWIDTH | OA_HEIGHT)
#define OA_PY_PWIDTH_PHEIGHT (OA_PY | OA_PWIDTH | OA_PHEIGHT)
#define OA_PX_PY (OA_PX | OA_PY)
#define OA_PX_PY_HEIGHT (OA_PX | OA_PY | OA_HEIGHT)
#define OA_PX_PY_PHEIGHT (OA_PX | OA_PY | OA_PHEIGHT)
#define OA_PX_PY_PWIDTH (OA_PX | OA_PY | OA_PWIDTH)
#define OA_PX_PY_PWIDTH_PHEIGHT (OA_PX | OA_PY | OA_PWIDTH | OA_PHEIGHT)
#define OA_PX_PY_WIDTH (OA_PX | OA_PY | OA_WIDTH)
#define OA_PX_PY_WIDTH_HEIGHT (OA_PX | OA_PY | OA_WIDTH | OA_HEIGHT)
#define OA_PX_Y (OA_PX | OA_Y)
#define OA_PX_Y_PWIDTH (OA_PX | OA_Y | OA_PWIDTH)
#define OA_PX_Y_PHEIGHT (OA_PX | OA_Y | OA_PHEIGHT)
#define OA_X_Y (OA_X | OA_Y)
#define OA_X_HEIGHT (OA_X | OA_HEIGHT)
#define OA_X_PHEIGHT (OA_X | OA_PHEIGHT)
#define OA_X_WIDTH (OA_X | OA_WIDTH)
#define OA_X_PWIDTH (OA_X | OA_PWIDTH)
#define OA_X_PY (OA_X | OA_PY)
#define OA_X_PY_PHEIGHT (OA_X | OA_PY | OA_PHEIGHT)
#define OA_Y_PWIDTH (OA_Y | OA_PWIDTH)
#define OA_Y_WIDTH (OA_Y | OA_WIDTH)
#define TRAY_ICON_MSG WM_APP + 1
//#define GCL_HBRBACKGROUND -10
#define CBXS_DISABLED 4l
#define CBXS_HOT 2l
#define CBXS_NORMAL 1l
#define CBXS_PRESSED 3l
#define CP_DROPDOWNBUTTON 1l
#define ETDT_DISABLE 0x01
#define ETDT_ENABLE 0x02
#define ETDT_ENABLETAB 0x06
#define ETDT_USETABTEXTURE 0x04
#define STAP_ALLOW_CONTROLS 0x02
#define STAP_ALLOW_NONCLIENT 0x01
#define STAP_ALLOW_WEBCONTENT 0x04
#define WM_THEMECHANGED 0x031A
