///////////////////////////////////////////////////////////////////////////
// Set.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET Set()-related preprocessor directives
//

#define _SET_EXACT        1
#define _SET_FIXED        2     // SetFixed()       LOGIC
#define _SET_DECIMALS     3     // SetDecimals()    INT
#define _SET_DATEFORMAT   4     // SetDateFormat()  STRING
#define _SET_EPOCH        5     // SetEpoch()       INT
#define _SET_PATH         6     // SetPath()        STRING
#define _SET_DEFAULT      7     // SetDefault()     STRING
#define _SET_EXCLUSIVE    8     // SetExclusive()   LOGIC
#define _SET_SOFTSEEK     9     // SetSoftseek()    LOGIC
#define _SET_UNIQUE      10     // SetUnique()      LOGIC
#define _SET_DELETED     11     // SetDeleted()     LOGIC
#define _SET_CANCEL      12     // SetCancel()      LOGIC
#define _SET_DEBUG       13
#define _SET_TYPEAHEAD   14     // SetTypeahead()   INT
#define _SET_COLOR       15     // SetColor()       STRING
#define _SET_CURSOR      16     // SetCursor()      INT
#define _SET_CONSOLE     17     // SetConsole()     LOGIC
#define _SET_ALTERNATE   18     // SetAlternate()   LOGIC
#define _SET_ALTFILE     19     // SetAltFile()     STRING
#define _SET_DEVICE      20     // SetDevice()      STRING
#define _SET_EXTRA       21     // SetExtra()       LOGIC
#define _SET_EXTRAFILE   22     // SetExtraFile()   STRING
#define _SET_PRINTER     23     // SetPrinter()     LOGIC
#define _SET_PRINTFILE   24     // SetPrintFile()   STRING
#define _SET_MARGIN      25     // SetMargin()      INT
#define _SET_BELL        26     // SetBell()        LOGIC
#define _SET_CONFIRM     27     // SetConfirm()     LOGIC
#define _SET_ESCAPE      28     // SetEscape()      LOGIC
#define _SET_INSERT      29     // SetInsert()      LOGIC
#define _SET_EXIT        30     // SetExit()        LOGIC
#define _SET_INTENSITY   31     // SetIntensity()   LOGIC
#define _SET_SCOREBOARD  32     // SetScoreboard()  LOGIC
#define _SET_DELIMITERS  33     // SetDelimiters()  STRING
#define _SET_DELIMCHARS  34     // SetDelimChars()  STRING
#define _SET_WRAP        35     // SetWrap()        LOGIC
#define _SET_MESSAGE     36     // SetMessage()     INT
#define _SET_MCENTER     37     // SetMCenter()     LOGIC
#define _SET_SCROLLBREAK 38     // SetScrollBreak() LOGIC
#define _SET_DIGITS      39     // SetDigits()      INT
#define _SET_NETERR      40
#define _SET_HPLOCK      41
// ??                    42
// ??                    43
#define _SET_ANSI        44
#define _SET_YIELD       45
#define _SET_LOCKTRIES   46     // LockTries()      INT
// ??                    47-97
#define _SET_DICT        98
#define _SET_INTL        99

#define _SET_COUNT       99


// eof
