///////////////////////////////////////////////////////////////////////////
// VOSystemClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// System Classes library
//

#define ccOptimistic 1
#define ccNone 0
#define ccStable 2
#define ccRepeatable 3
#define ccFile 4
#define ccUser 1000
#define DBC_INDEXNAME 1
#define DBC_INDEXPATH 2
#define DBC_ORDERS 3
#define DBC_TAGNAME 1
#define DBC_DUPLICATE 2
#define DBC_ASCENDING 3
#define DBC_KEYEXP 4
#define DBC_FOREXP 5
#define DBC_SYMBOL 1
#define DBC_NAME 2
#define DBC_FIELDSPEC 3
#define NOTIFYFIELDCHANGE -1
#define NOTIFYCLEARRELATION 25
#define NOTIFYCLOSE 0
#define NOTIFYCOMPLETION 1
#define NOTIFYINTENTTOMOVE 2
#define NOTIFYRECORDCHANGE 3
#define NOTIFYGOBOTTOM 4
#define NOTIFYGOTOP 5
#define NOTIFYDELETE 6
#define NOTIFYAPPEND 7
#define NOTIFYFILECHANGE 10
#define NOTIFYRELATIONCHANGE 20
#define NOTIFYCONCURRENCYCONTROLMODE 50
#define TYPE_MULTIMEDIA 42
#ifndef MAXFILENAME
   #define MAXFILENAME 260
#endif
#define MAXEXTNAME 128
#define MAXDIRNAME 256
#define MAXDRIVENAME 128
