#ifndef GlobalDefines

#define GlobalDefines

#DEFINE WIN32SUCCESS 0

#define AEF_REC_APPBODY 0x010F
#define AEF_REC_APPDESC 0x000F
#define AEF_REC_APPEXPNAME 0x0126
#define AEF_REC_APPNAME 0x0002
#define AEF_REC_CH 0x0125
#define AEF_REC_CHFILE 0x0124
#define AEF_REC_DLL (0x0060 )
#define AEF_REC_DLLFILE 0x0102
#define AEF_REC_DLLFLG 0x000B
#define AEF_REC_END 0xffff
#define AEF_REC_ENTBODY 0x010D
#define AEF_REC_ENTNAME 0x0040
#define AEF_REC_EXENAME 0x000D
#define AEF_REC_EXTMOD 0x0101
#define AEF_REC_EXTMODNAME 0x0022
#define AEF_REC_EXTRES (0x0103 )
#define AEF_REC_EXTRESNAME 0x0061
#define AEF_REC_GROUPNAME 0x0108
#define AEF_REC_HEADER 1
#define AEF_REC_LIBFLG 0x000A
#define AEF_REC_MODBODY 0x010E
#define AEF_REC_MODEXPNAME 0x0127
#define AEF_REC_MODNAME 0x0020
#define AEF_REC_SPATH 0x0004
#define AEF_REC_UDC 0x0005
#define AEF_REC_UDCFILE (0x0100 )

#define FabAEFFileFILE_TEXT "CA-VO Application Export File"
#define FabAEFFileFILE_TEXT_LEN 30
#define FabAEFFileFILE_VERSION_10 (_CHR(0)+_CHR(1))
#define FabAEFFileFILE_VERSION_20 (_CHR(0)+_CHR(2))
#define FabAEFFileFILE_VERSION_LEN 2
#define FabFabAEFFileFile_REC_TIME (0x0006 )

#define MEFFILE_TEXT "CA-VO Module Export File"
#define MEFFILE_TEXT_LEN 25
#define MEFFILE_VERSION_10 FabAEFFileFILE_VERSION_10
#define MEFFILE_VERSION_20 FabAEFFileFILE_VERSION_20
#define MEFFILE_VERSION_LEN 2
#define MEF_ENT_CREATETIME 5
#define MEF_ENT_LASTBUILD 4
#define MEF_ENT_NAME 1
#define MEF_ENT_PROTO 3
#define MEF_ENT_PTR 2
#define MEF_ENT_SIZE 5
#define MEF_REC_ENTPROTO 0x004e
#define MEF_REC_ENTSOURCE 0x0041


#endif
