///////////////////////////////////////////////////////////////////////////
// VOReportClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// Report Classes library
//

#define WRM_NTFY_MSG_BASE 6500
#define MAX_RCC_FONT 2
#define MAX_RCC_COLOR 12
#define CAWRM_NTFY_CLOSE (WM_USER+1)
#define CAWRM_NTFY_NEW_WRAP (WM_USER+2)
#define CAWRM_NTFY_COMMAND (WM_USER+3)
#define CAWRM_NTFY_SET_MENU (WM_USER+4)
#define CAWRM_NTFY_ADVISE (WM_USER+5)
#define CAWRM_NTFY_DEPENDENCY (WM_USER+6)
#define CAWRM_NTFY_PREVIEW (WM_USER+7)
#define CAWRM_NTFY_ADVISE_CLEAR (WM_USER+9)
#define CAWRM_NTFY_ABOUT (WM_USER+10)
#define CAWRM_NTFY_EDIT_QUERY (WM_USER+8)
#define CAWRM_NTFY_HELP (WM_USER+11)
#define CAWRM_NTFY_SAVE (WM_USER+12)
#define WRM_NTFY_ADVISE_CLEAR (WRM_NTFY_MSG_BASE+CAWRM_NTFY_ADVISE_CLEAR)
#define TP_MENU_BASE 100
#define NTFY_MSG_BASE 2000
#define DBA_MENU_BASE (TP_MENU_BASE +1600)
#define QQ_MENU_BASE (TP_MENU_BASE +400)
#define RET_REPORT_OPEN 1
#define RET_FILE_NAME 1
#define CAWRMWRAPINFO_WRMTYPE 2
#define REPORTCLOSEEVENT 301
#define REPORTCOMPLETEERROREVENT 305
#define REPORTCOMPLETEEVENT 302
#define REPORTFILESAVEEVENT 306
#define REPORTOPENEVENT 300
#define REPORTSERVERCLOSEEVENT 303
#define REPORTVIEWCLOSEEVENT 304
#define RET_RPTEVT_REPORT_OPENED 1
#define RET_RPTEVT_PRINTER_CANCELED 2
#define RET_RPTEVT_REPORT_COMPLETE 3
#define RET_RPTEVT_REPORT_CLOSE 4
#define RET_RPTEVT_FILE_SAVE 5
#define RET_RPTEVT_VIEW_CLOSE 6
#define RET_REPORT_CREATE 0
#define RPTSTYLE_TABULAR 2
#define RET_QUERY_CQMSQLSTRING 4
#define RPTSTYLE_FREESTYLE 1
#define RPTSTYLE_FORM 3
#define RPTSTYLE_LABEL 4
#define RPTSTYLE_LETTER 5
#define RPTSTYLE_CROSSTAB 6
#define RPTSTYLE_NOTSPECIFIED 0
#define FILE_NEW 1
#define FILE_OPEN 2
#define WRM_NTFY_CLOSE (WRM_NTFY_MSG_BASE+CAWRM_NTFY_CLOSE)
#define WRM_NTFY_NEW_WRAP (WRM_NTFY_MSG_BASE+CAWRM_NTFY_NEW_WRAP)
#define WRM_NTFY_COMMAND (WRM_NTFY_MSG_BASE+CAWRM_NTFY_COMMAND)
#define WRM_NTFY_SET_MENU (WRM_NTFY_MSG_BASE+CAWRM_NTFY_SET_MENU)
#define WRM_NTFY_ADVISE (WRM_NTFY_MSG_BASE+CAWRM_NTFY_ADVISE)
#define WRM_NTFY_DEPENDENCY (WRM_NTFY_MSG_BASE+CAWRM_NTFY_DEPENDENCY)
#define WRM_NTFY_PREVIEW (WRM_NTFY_MSG_BASE+CAWRM_NTFY_PREVIEW)
#define WRM_NTFY_EDIT_QUERY (WRM_NTFY_MSG_BASE+CAWRM_NTFY_EDIT_QUERY)
#define WRM_NTFY_ABOUT (WRM_NTFY_MSG_BASE +CAWRM_NTFY_ABOUT)
#define WRM_NTFY_HELP (WRM_NTFY_MSG_BASE +CAWRM_NTFY_HELP)
#define WRM_NTFY_SAVE (WRM_NTFY_MSG_BASE +CAWRM_NTFY_SAVE)
