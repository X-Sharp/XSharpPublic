#define DIR_HREF_STOP ">"
///////////////////////////////////////////////////////////////////////////
// VOInternetClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// Internet Classes library
//

#define HEADER_ACCEPT "Accept: *" + "/" + "*" + CRLF + CRLF
#define HEADER_ACCEPT_REQ "*" + "/" + "*"
#define URL_LOCAL_HOST "http://localhost"
#define DIR_HREF_START "<A HREF="
#define TEMP_MESSAGES "MESSAGES"
#define TEMP_RFC_SIZE "(RFC822.SIZE"
#define NOTIFY_CINetDial_ERROR 1
#define NOTIFY_CINetDial_QueryHangUp 2
#define NOTIFY_CINetDial_CONNECTED 3
#define NOTIFY_CINetDial_DISCONNECTED 4
#define NOTIFY_CINetDial_QueryHangUpAll 5
#define NEWSLIST_FIRST 3
#define NEWSLIST_LAST 2
#define NEWSLIST_MAX 4
#define NEWSLIST_NAME 1
#define NEWSLIST_POST 4
#define STATUS_HANDLE 1
#define STATUS_OP 2
#define STATUS_SIZE 1024
#define FIOASYNC 0x8004667D
#define FIONBIO 0x8004667E
#define FIONREAD 0x4004667F
#define INVALID_SOCKET 0xFFFFFFFFU
#define MIN_SOCKETS_REQUIRED 10
#define SCMD_NEWSOCKETACCEPTED -101
#define SCMD_SOCKETSTATUSCHANGED -100
#define SD_BOTH 2
#define SD_RECEIVE 0
#define SD_SEND 1
#define SOCK_BLOCK_SIZE 520
#define SSTAT_CONNECTED 5
#define SSTAT_CONNECTING 2
#define SSTAT_DISCONNECTED 1
#define SSTAT_DISCONNECTING 4
#define SSTAT_ERRORSTATE 6
#define SSTAT_LISTENING 3
#define SSTAT_TIMEDOUT 7
#define SSTAT_UNINITIALIZED 0
#define WS_VERSION_MAJOR 1
#define WS_VERSION_MINOR 1
#define WS_VERSION_REQUIRED 0x0101
#define ATTACHID_PATHFLAG ">"
#define ATTACH_BEGIN BOUNDARY_DELIMITER
#define ATTACH_CONTENTID 2
#define ATTACH_CONTENTTYPE 5
#define ATTACH_FILENAME 4
#define ATTACH_FILESIZE 3
#define ATTACH_FULLPATH 7
#define ATTACH_SIZE 8
#define ATTACH_STOREID 1
#define ATTACH_TRANSFERENCODING 6
#define ATTACHMENT_END BOUNDARY_DELIMITER + CRLF + CRLF + "." + CRLF
#define BOUNDARY_DELIMITER "--"
#define BOUNDARY_START CRLF + BOUNDARY_DELIMITER
#define BOUNDARY_VO_ID "Visual_Objects_BOUNDARY"
#define BOUNDARY_VO "===" + BOUNDARY_VO_ID + "==="
#define BOUNDARY_VO_ID "Visual_Objects_BOUNDARY"
#define CHARSET_ISO "iso-8859-"
#define CHARSET_ISO1 e"\"" + CHARSET_ISO + e"1\""
#define CHARSET_USASCII "us-ascii"
#define CHARSET_UTF8 "utf-8"
#define CLOSING_CONNECTION 4
#define CODING_7BIT "7bit"
#define CODING_8BIT "8bit"
#define CODING_BASE64 "base64"
#define CODING_QP "quoted-printable"
#define CODING_TYPE_7BIT 4
#define CODING_TYPE_8BIT 5
#define CODING_TYPE_BASE64 2
#define CODING_TYPE_NONE 0
#define CODING_TYPE_PRINTABLE 3
#define CODING_TYPE_UNKNOWN 5
#define CODING_TYPE_UUENCODE 1
#define CODING_UUENCODE "uuencode"
#define CONNECTED 12
#define CONNECTING 1
#define CONTENT_APPLICATION "application/octet-stream"
#define CONTENT_AUDIO "audio"
#define CONTENT_DEFAULT "text/plain; charset=us-ascii"
#define CONTENT_IMAGE "image"
#define CONTENT_MESSAGE "message"
#define CONTENT_MULTIPART "multipart"
#define CONTENT_MULTIPART_ALTERNATE CONTENT_MULTIPART + "/alternative"
#define CONTENT_MULTIPART_MIXED CONTENT_MULTIPART + "/mixed"
#define CONTENT_MULTIPART_RELATED CONTENT_MULTIPART + "/related"
#define CONTENT_MULTIPART_REPORT CONTENT_MULTIPART + "/report"
#define CONTENT_TEXT "text"
#define CONTENT_TEXT_HTML CONTENT_TEXT + "/html"
#define CONTENT_TEXT_PLAIN CONTENT_TEXT+"/plain"
#define CONTENT_VIDEO "video"
#define DEFAULT_BOUNDARY CRLF + CRLF
#define DEFAULT_STOPDATA CRLF + "." + CRLF
#define EMAIL_FORMAT_MIME 2
#define EMAIL_FORMAT_UUENCODE 1
#define ERR_FILE_EXISTS INTERNET_ERROR_BASE + 224
#define ERR_LOGON_FAILED INTERNET_ERROR_BASE + 223
#define ERR_NEWSGROUP_MISSING INTERNET_ERROR_BASE + 411
#define ERR_NO_ARTICLE INTERNET_ERROR_BASE + 430
#define ERR_NO_ARTICLE_NUMBER INTERNET_ERROR_BASE + 423
#define ERR_NO_ARTICLE_SELECTED INTERNET_ERROR_BASE + 420
#define ERR_NO_NEWSGROUP INTERNET_ERROR_BASE + 412
#define ERR_UNKNOWN_CODE_TYPE INTERNET_ERROR_BASE + 225
#define ERR_WSA_WAIT_TIMEOUT 12258
#define ESTABLISHING_SESSION 2
#define IMAGE_BMP "image/bmp"
#define IMAGE_JPEG "image/jpeg"
#define IMAGE_JPG "image/jpg"
#define IMAGE_TYPE "image"
#define IPPORT_IMAP 143
#define IPPORT_NNTP 119
#define IPPORT_POP 110
#define LOGGED_OFF 11
#define LOGGED_ON 10
#define LOGGING_ON 6
#define MAX_SOCKBUFF 2500
#define MIME_MULTI_PART "This is a multi-part message in MIME format."
#define MY_STOPDATA CRLF + ".." +CRLF
#define RETREIVING_DATA 8
#define SENDING_DATA 9
#define SENDING_HEADER 3
#define SENDING_REQUEST 7
#define TAB _CHR(9)
#define TEMP_ATTACHMENT "attachment"
#define TEMP_BCC "Bcc:"
#define TEMP_BOUNDARY "boundary="
#define TEMP_BOUND TEMP_BOUNDARY + e"\""
#define TEMP_CC "Cc:"
#define TEMP_CHARSET "charset="
#define TEMP_CONTENT "Content-Type:"
#define TEMP_CONTENTDISPOSITION "Content-Disposition:"
#define TEMP_CONTENTID "Content-Id:"
#define TEMP_DATE "Date:"
#define TEMP_DECODE_BOUND CRLF+CRLF
#define TEMP_DISPOSITIONNOTIFICATION "Disposition-Notification-To:"
#define TEMP_ENCODE "Content-Transfer-Encoding:"
#define TEMP_FNAME "filename="
#define TEMP_FOLLOWUP "Followup-To:"
#define TEMP_FROM "From:"
#define TEMP_MAILER "X-Mailer:"
#define TEMP_MESSAGEID "Message-ID:"
#define TEMP_MIMEVERSION "Mime-Version: 1.0"
#define TEMP_MULIPARTINFO "This is a multi-part message in MIME format."
#define TEMP_NAME "name="
#define TEMP_NEWSGROUPS "Newsgroups:"
#define TEMP_ORGANIZATION "Organization:"
#define TEMP_PATH "Path:"
#define TEMP_POSTED "Posted:"
#define TEMP_PRIORITY "X-Priority:"
#define TEMP_REFERENCES "References:"
#define TEMP_REPLY "Reply-To:"
#define TEMP_RETURN_RECEIPT "Return-Receipt-To:"
#define TEMP_SENDER "Sender:"
#define TEMP_STOP e"\""
#define TEMP_SUBJECT "Subject:"
#define TEMP_TO "To:"
#define UUE_END CRLF + "end"
#define UUE_START_EMAIL "begin 777 "
#define UUE_START_NEWS "begin"
#define UUE_STOP _CHR(96) + CRLF
#define WAITING_FOR_ACTION 5
#define WSA_WAIT_TIMEOUT STATUS_TIMEOUT
#define WSABASEERR 10000
#define WSAEACCES WSABASEERR+13
#define WSAEADDRINUSE WSABASEERR+48
#define WSAEADDRNOTAVAIL WSABASEERR+49
#define WSAEAFNOSUPPORT WSABASEERR+47
#define WSAEALREADY WSABASEERR+37
#define WSAEBADF WSABASEERR+9
#define WSAECONNABORTED WSABASEERR+53
#define WSAECONNREFUSED WSABASEERR+61
#define WSAECONNRESET WSABASEERR+54
#define WSAEDESTADDRREQ WSABASEERR+39
#define WSAEDISCON WSABASEERR+101
#define WSAEDQUOT WSABASEERR+69
#define WSAEFAULT WSABASEERR+14
#define WSAEHOSTDOWN WSABASEERR+64
#define WSAEHOSTUNREACH WSABASEERR+65
#define WSAEINPROGRESS WSABASEERR+36
#define WSAEINTR WSABASEERR+4
#define WSAEINVAL WSABASEERR+22
#define WSAEISCONN WSABASEERR+56
#define WSAELOOP WSABASEERR+62
#define WSAEMFILE WSABASEERR+24
#define WSAEMSGSIZE WSABASEERR+40
#define WSAENAMETOOLONG WSABASEERR+63
#define WSAENETDOWN WSABASEERR+50
#define WSAENETRESET WSABASEERR+52
#define WSAENETUNREACH WSABASEERR+51
#define WSAENOBUFS WSABASEERR+55
#define WSAENOPROTOOPT WSABASEERR+42
#define WSAENOTCONN WSABASEERR+57
#define WSAENOTEMPTY WSABASEERR+66
#define WSAENOTSOCK WSABASEERR+38
#define WSAEOPNOTSUPP WSABASEERR+45
#define WSAEPFNOSUPPORT WSABASEERR+46
#define WSAEPROCLIM WSABASEERR+67
#define WSAEPROTONOSUPPORT WSABASEERR+43
#define WSAEPROTOTYPE WSABASEERR+41
#define WSAEREMOTE WSABASEERR+71
#define WSAESHUTDOWN WSABASEERR+58
#define WSAESOCKTNOSUPPORT WSABASEERR+44
#define WSAESTALE WSABASEERR+70
#define WSAETIMEDOUT WSABASEERR+60
#define WSAETOOMANYREFS WSABASEERR+59
#define WSAEUSERS WSABASEERR+68
#define WSAEWOULDBLOCK WSABASEERR+35
#define WSAHOST_NOT_FOUND WSABASEERR+1001
#define WSANO_DATA WSABASEERR+1004
#define WSANO_ADDRESS WSANO_DATA
#define WSANO_RECOVERY WSABASEERR+1003
#define WSANOTINITIALISED WSABASEERR+93
#define WSASYSNOTREADY WSABASEERR+91
#define WSATRY_AGAIN WSABASEERR+1002
#define WSAVERNOTSUPPORTED WSABASEERR+92
