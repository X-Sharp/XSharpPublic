///////////////////////////////////////////////////////////////////////////
// VOWin32APILibrary.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// Windows API library
//

#define CTS_READONLY 0x00000100
#define CTS_SINGLESEL 0x00000200
#define CTS_MULTIPLESEL 0x00000400
#define CTS_EXTENDEDSEL 0x00000800
#define CTS_BLOCKSEL 0x00001000
#define CTS_SPLITBAR 0x00002000
#define CTS_VERTSCROLL 0x00004000
#define CTS_HORZSCROLL 0x00008000
#define CTS_INTEGRALWIDTH 0x00000001
#define CTS_INTEGRALHEIGHT 0x00000002
#define CTS_EXPANDLASTFLD 0x00000004
#define CTS_ASYNCNOTIFY 0x00000080
#define CN_ASSOCIATEGAIN 501
#define CN_ASSOCIATELOSS 502
#define CN_RANGECHANGE 503
#define CN_BEGTTLEDIT 504
#define CN_ENDTTLEDIT 505
#define CN_BEGFLDTTLEDIT 506
#define CN_ENDFLDTTLEDIT 507
#define CN_BEGRECEDIT 508
#define CN_ENDRECEDIT 509
#define CN_BEGFLDEDIT 510
#define CN_ENDFLDEDIT 511
#define CN_EMPHASIS 512
#define CN_SETFOCUS 513
#define CN_KILLFOCUS 514
#define CN_QUERYDELTA 515
#define CN_ENTER 516
#define CN_INSERT 517
#define CN_DELETE 518
#define CN_ESCAPE 519
#define CN_TAB 520
#define CN_RECSELECTED 521
#define CN_RECUNSELECTED 522
#define CN_CHARHIT 523
#define CN_ROTTLDBLCLK 524
#define CN_ROFLDTTLDBLCLK 525
#define CN_ROFLDDBLCLK 526
#define CN_NEWFOCUS 527
#define CN_NEWFOCUSREC 528
#define CN_NEWFOCUSFLD 529
#define CN_QUERYFOCUS 530
#define CN_F1 531
#define CN_F2 532
#define CN_F3 533
#define CN_F4 534
#define CN_F5 535
#define CN_F6 536
#define CN_F7 537
#define CN_F8 538
#define CN_F9 539
#define CN_F10 540
#define CN_F11 541
#define CN_F12 542
#define CN_F13 543
#define CN_F14 544
#define CN_F15 545
#define CN_F16 546
#define CN_F17 547
#define CN_F18 548
#define CN_F19 549
#define CN_F20 550
#define CN_F21 551
#define CN_F22 552
#define CN_F23 553
#define CN_F24 554
#define CN_TTLBTNCLK 555
#define CN_FLDTTLBTNCLK 556
#define CN_VSCROLL_TOP 557
#define CN_VSCROLL_BOTTOM 558
#define CN_VSCROLL_PAGEUP 559
#define CN_VSCROLL_PAGEDOWN 560
#define CN_VSCROLL_LINEUP 561
#define CN_VSCROLL_LINEDOWN 562
#define CN_VSCROLL_THUMBPOS 563
#define CN_HSCROLL_PAGEUP 564
#define CN_HSCROLL_PAGEDOWN 565
#define CN_HSCROLL_LINEUP 566
#define CN_HSCROLL_LINEDOWN 567
#define CN_HSCROLL_THUMBPOS 568
#define CN_FLDSIZED 569
#define CN_FLDMOVED 570
#define CN_FLDSELECTED 571
#define CN_FLDUNSELECTED 572
#define CN_SPLITBAR_CREATED 573
#define CN_SPLITBAR_MOVED 574
#define CN_SPLITBAR_DELETED 575
#define CN_NEWRECSELECTLIST 576
#define CN_BGNRECSELECTION 577
#define CN_ENDRECSELECTION 578
#define CN_NEWFLDSELECTLIST 579
#define CN_BGNFLDSELECTION 580
#define CN_ENDFLDSELECTION 581
#define CN_LK_ARROW_UP 582
#define CN_LK_ARROW_DOWN 583
#define CN_LK_ARROW_LEFT 584
#define CN_LK_ARROW_RIGHT 585
#define CN_LK_HOME 586
#define CN_LK_END 587
#define CN_LK_PAGEUP 588
#define CN_LK_PAGEDOWN 589
#define CN_LK_NEWFOCUS 590
#define CN_LK_NEWFOCUSREC 591
#define CN_LK_NEWFOCUSFLD 592
#define CN_LK_VS_TOP 593
#define CN_LK_VS_BOTTOM 594
#define CN_LK_VS_PAGEUP 595
#define CN_LK_VS_PAGEDOWN 596
#define CN_LK_VS_LINEUP 597
#define CN_LK_VS_LINEDOWN 598
#define CN_LK_VS_THUMBPOS 599
#define CN_LK_HS_PAGEUP 600
#define CN_LK_HS_PAGEDOWN 601
#define CN_LK_HS_LINEUP 602
#define CN_LK_HS_LINEDOWN 603
#define CN_LK_HS_THUMBPOS 604
#define CN_OWNERSETFOCUSTOP 605
#define CN_OWNERSETFOCUSBOT 606
#define CN_CUT 607
#define CN_COPY 608
#define CN_PASTE 609
#define CN_CLEAR 610
#define CN_UNDO 611
#define CN_RBTNCLK 612
#define CN_VSCROLL_THUMBTRK 613
#define CN_FLDSIZECHANGED 614
#define CN_SIZECHANGED 615
#define LAST_CN_MSG 3000
#define CNTCOLOR_TITLE 0
#define CNTCOLOR_FLDTITLES 1
#define CNTCOLOR_TEXT 2
#define CNTCOLOR_GRID 3
#define CNTCOLOR_CNTBKGD 4
#define CNTCOLOR_HIGHLIGHT 5
#define CNTCOLOR_HITEXT 6
#define CNTCOLOR_TTLBKGD 7
#define CNTCOLOR_FLDTTLBKGD 8
#define CNTCOLOR_FLDBKGD 9
#define CNTCOLOR_3DHIGH 10
#define CNTCOLOR_3DSHADOW 11
#define CNTCOLOR_TTLBTNTXT 12
#define CNTCOLOR_TTLBTNBKGD 13
#define CNTCOLOR_FLDBTNTXT 14
#define CNTCOLOR_FLDBTNBKGD 15
#define CNTCOLOR_UNUSEDBKGD 16
#define CNTCOLOR_INUSE 17
#define CNTCOLORS 18
#define CF_GENERAL 0
#define CF_TITLE 1
#define CF_FLDTITLE 2
#define CC_GENERAL 0
#define CC_TITLE 1
#define CC_FLDTITLE 2
#define CFM_LEFT 0
#define CFM_RIGHT 1
#define CFM_UP 2
#define CFM_DOWN 3
#define CFM_PAGEUP 4
#define CFM_PAGEDOWN 5
#define CFM_FIRSTFLD 6
#define CFM_LASTFLD 7
#define CFM_HOME 8
#define CFM_END 9
#define CFM_NEXTSPLITWND 10
#define CB_LEFT 0
#define CB_RIGHT 1
#define AS_AVGCHAR 1
#define AS_MAXCHAR 2
#define AS_PIXELS 3
#define BK_GENERAL 0
#define BK_UNUSED 1
#define BK_TITLE 2
#define BK_FLDTITLE 3
#define BK_FLD 4
#define CSB_SHOW 0
#define CSB_LEFT 1
#define CSB_MIDDLE 2
#define CSB_RIGHT 3
#define CSB_XCOORD 4
#define CSB_FIRST 5
#define CSB_LAST 6
#define CSB_NEXT 7
#define CSB_PREV 8
#define CA_LS_NONE 0
#define CA_LS_NARROW 1
#define CA_LS_MEDIUM 2
#define CA_LS_WIDE 3
#define CA_LS_DOUBLE 4
#define CE_ID_EDIT1 1001
#define CE_ID_EDIT2 1002
#define CE_ID_EDIT3 1003
#define CE_ID_EDIT4 1004
#define CE_ID_EDIT5 1005
#define CE_ID_EDIT6 1006
#define CE_ID_EDIT7 1007
#define CE_ID_EDIT8 1008
#define CE_ID_EDIT9 1009
#define CE_ID_EDIT10 1010
#define CE_ID_EDIT11 1011
#define CE_ID_EDIT12 1012
#define CV_ICON 0x0001
#define CV_NAME 0x0002
#define CV_TEXT 0x0004
#define CV_DETAIL 0x0008
#define CV_MINI 0x0010
#define CV_FLOW 0x0020
#define CA_TA_TOP 0x00000001
#define CA_TA_VCENTER 0x00000002
#define CA_TA_BOTTOM 0x00000004
#define CA_TA_LEFT 0x00000008
#define CA_TA_HCENTER 0x00000010
#define CA_TA_RIGHT 0x00000020
#define CA_TTLREADONLY 0x00000001
#define CA_TITLE 0x00000002
#define CA_FLDTITLES 0x00000004
#define CA_OWNERPNTBK 0x00000008
#define CA_OWNERPNTUNBK 0x00000010
#define CA_TTLSEPARATOR 0x00000020
#define CA_FLDSEPARATOR 0x00000040
#define CA_RECSEPARATOR 0x00000080
#define CA_DRAWBMP 0x00000100
#define CA_DRAWICON 0x00000200
#define CA_TTLBTNPRESSED 0x00000400
#define CA_TITLE3D 0x00000800
#define CA_FLDTTL3D 0x00001000
#define CA_VERTFLDSEP 0x00002000
#define CA_TRANTTLBMP 0x00004000
#define CA_TRANTTLBTNBMP 0x00008000
#define CA_OWNERVSCROLL 0x00010000
#define CA_SIZEABLEFLDS 0x00020000
#define CA_MOVEABLEFLDS 0x00040000
#define CA_APPSPLITABLE 0x00080000
#define CA_OWNERPNTTTLBK 0x00100000
#define CA_WIDEFOCUSRECT 0x00200000
#define CA_HSCROLLBYCHAR 0x00400000
#define CA_WANTVTHUMBTRK 0x00800000
#define CA_DYNAMICVSCROLL 0x01000000
#define CFA_FLDREADONLY 0x00000001
#define CFA_FLDTTLREADONLY 0x00000002
#define CFA_HORZSEPARATOR 0x00000004
#define CFA_VERTSEPARATOR 0x00000008
#define CFA_CURSORED 0x00000010
#define CFA_FLDTTL3D 0x00000020
#define CFA_TRANFLDTTLBMP 0x00000040
#define CFA_OWNERDRAW 0x00000080
#define CFA_HEX 0x00000100
#define CFA_OCTAL 0x00000200
#define CFA_BINARY 0x00000400
#define CFA_SCIENTIFIC 0x00000800
#define CFA_TRANFLDBTNBMP 0x00001000
#define CFA_FLDBTNPRESSED 0x00002000
#define CFA_SIZEABLEFLD 0x00004000
#define CFA_MOVEABLEFLD 0x00008000
#define CFA_NONSIZEABLEFLD 0x00010000
#define CFA_NONMOVEABLEFLD 0x00020000
#define CFA_OWNERPNTFTBK 0x00040000
#define CFA_OWNERPNTFLDBK 0x00080000
#define CFT_STRING 0
#define CFT_LPSTRING 1
#define CFT_WORD 2
#define CFT_UINT 3
#define CFT_INT 4
#define CFT_DWORD 5
#define CFT_LONG 6
#define CFT_FLOAT 7
#define CFT_DOUBLE 8
#define CFT_BCD 9
#define CFT_DATE 10
#define CFT_TIME 11
#define CFT_BMP 12
#define CFT_ICON 13
#define CFT_CAMASK 14
#define CFT_CANUMBER 15
#define CFT_CADATE 16
#define CFT_CATIME 17
#define CFT_CUSTOM 18
#define CFT_CHAR 19
#define CFT_CANUMBERUNSGN 20
#define CRA_RECREADONLY 0x00000001
#define CRA_CURSORED 0x00000002
#define CRA_DROPONABLE 0x00000004
#define CRA_FILTERED 0x00000008
#define CRA_FLDSELECTED 0x00000010
#define CRA_SELECTED 0x00000020
#define CRA_TARGET 0x00000040
#define CRA_FIRSTREC 0x00000080
#define CRA_LASTREC 0x00000100
#define CRA_INUSE 0x00000200
#define MAX_BTNTXT_LEN 64
#define MAX_SPLITBARS 20
#define CASPLIT_CLASS "CA_SplitWindow32"
#define SWS_HALIGN 0x00000001
#define SWS_VALIGN 0x00000002
#define SWS_TEXTHASPARMS 0x00000004
#define SWS_NOHORZDRAG 0x00000008
#define SWS_NOVERTDRAG 0x00000010
#define SWN_ASSOCIATEGAIN 401
#define SWN_ASSOCIATELOSS 402
#define SPLTCOLOR_BAR 0
#define SPLTCOLOR_BARFRAME 1
#define SPLTCOLOR_WINDOW 2
#define SPLTCOLOR_3DHIGH 3
#define SPLTCOLOR_3DSHADOW 4
#define SPS_SHOWPANE 1
#define SPS_HIDEPANE 2
#define SPS_SHOWROW 3
#define SPS_HIDEROW 4
#define SPS_SHOWCOLUMN 5
#define SPS_HIDECOLUMN 6
#define SPS_SHOWALLPANES 7
#define SPS_HIDEALLPANES 8
#define CDERR_DIALOGFAILURE 0xFFFF
#define CDERR_GENERALCODES 0x0000
#define CDERR_STRUCTSIZE 0x0001
#define CDERR_INITIALIZATION 0x0002
#define CDERR_NOTEMPLATE 0x0003
#define CDERR_NOHINSTANCE 0x0004
#define CDERR_LOADSTRFAILURE 0x0005
#define CDERR_FINDRESFAILURE 0x0006
#define CDERR_LOADRESFAILURE 0x0007
#define CDERR_LOCKRESFAILURE 0x0008
#define CDERR_MEMALLOCFAILURE 0x0009
#define CDERR_MEMLOCKFAILURE 0x000A
#define CDERR_NOHOOK 0x000B
#define CDERR_REGISTERMSGFAIL 0x000C
#define PDERR_PRINTERCODES 0x1000
#define PDERR_SETUPFAILURE 0x1001
#define PDERR_PARSEFAILURE 0x1002
#define PDERR_RETDEFFAILURE 0x1003
#define PDERR_LOADDRVFAILURE 0x1004
#define PDERR_GETDEVMODEFAIL 0x1005
#define PDERR_INITFAILURE 0x1006
#define PDERR_NODEVICES 0x1007
#define PDERR_NODEFAULTPRN 0x1008
#define PDERR_DNDMMISMATCH 0x1009
#define PDERR_CREATEICFAILURE 0x100A
#define PDERR_PRINTERNOTFOUND 0x100B
#define PDERR_DEFAULTDIFFERENT 0x100C
#define CFERR_CHOOSEFONTCODES 0x2000
#define CFERR_NOFONTS 0x2001
#define CFERR_MAXLESSTHANMIN 0x2002
#define FNERR_FILENAMECODES 0x3000
#define FNERR_SUBCLASSFAILURE 0x3001
#define FNERR_INVALIDFILENAME 0x3002
#define FNERR_BUFFERTOOSMALL 0x3003
#define FRERR_FINDREPLACECODES 0x4000
#define FRERR_BUFFERLENGTHZERO 0x4001
#define CCERR_CHOOSECOLORCODES 0x5000
#define TYMED_HGLOBAL 1
#define TYMED_FILE 2
#define TYMED_ISTREAM 4
#define TYMED_ISTORAGE 8
#define TYMED_GDI 16
#define TYMED_MFPICT 32
#define TYMED_ENHMF 64
#define TYMED_NULL 0
#define DATADIR_GET 1
#define DATADIR_SET 2
#define DROPEFFECT_NONE 0
#define DROPEFFECT_COPY 1
#define DROPEFFECT_MOVE 2
#define DROPEFFECT_LINK 4
#define DROPEFFECT_SCROLL 0x80000000
#define OLEMISC_RECOMPOSEONRESIZE 0x1
#define OLEMISC_ONLYICONIC 0x2
#define OLEMISC_INSERTNOTREPLACE 0x4
#define OLEMISC_STATIC 0x8
#define OLEMISC_CANTLINKINSIDE 0x10
#define OLEMISC_CANLINKBYOLE1 0x20
#define OLEMISC_ISLINKOBJECT 0x40
#define OLEMISC_INSIDEOUT 0x80
#define OLEMISC_ACTIVATEWHENVISIBLE 0x100
#define OLEMISC_RENDERINGISDEVICEINDEPENDENT 0x200
#define OLEMISC_INVISIBLEATRUNTIME 0x400
#define OLEMISC_ALWAYSRUN 0x800
#define OLEMISC_ACTSLIKEBUTTON 0x1000
#define OLEMISC_ACTSLIKELABEL 0x2000
#define OLEMISC_NOUIACTIVATE 0x4000
#define OLEMISC_ALIGNABLE 0x8000
#define OLEMISC_SIMPLEFRAME 0x10000
#define OLEMISC_SETCLIENTSITEFIRST 0x20000
#define OLEMISC_IMEMODE 0x40000
#define OLEMISC_IGNOREACTIVATEWHENVISIBLE 0x80000
#define OLEMISC_WANTSTOMENUMERGE 0x100000
#define OLEMISC_SUPPORTSMULTILEVELUNDO 0x200000
#define OLEGETMONIKER_ONLYIFTHERE 1
#define OLEGETMONIKER_FORCEASSIGN 2
#define OLEGETMONIKER_UNASSIGN 3
#define OLEGETMONIKER_TEMPFORUSER 4
#define OLEWHICHMK_CONTAINER 1
#define OLEWHICHMK_OBJREL 2
#define OLEWHICHMK_OBJFULL 3
#define PSSTATE_UNINIT 1
#define PSSTATE_SCRIBBLE 2
#define PSSTATE_HANDSOFF 3
#define STREAM_SEEK_SET 0
#define STREAM_SEEK_CUR 1
#define STREAM_SEEK_END 2
#define PSSTATE_ZOMBIE 4
#define OLERENDER_NONE 0
#define OLERENDER_DRAW 1
#define OLERENDER_FORMAT 2
#define OLERENDER_ASIS 3
#define ADVF_NODATA 1
#define ADVF_PRIMEFIRST 2
#define ADVF_ONLYONCE 4
#define ADVF_DATAONSTOP 64
#define ADVFCACHE_NOHANDLER 8
#define ADVFCACHE_FORCEBUILTIN 16
#define ADVFCACHE_ONSAVE 32
#define CLSCTX_REMOTE_SERVER 16
#define CLSCTX_INPROC_SERVER 1
#define CLSCTX_LOCAL_SERVER 4
#define CLSCTX_SERVER (CLSCTX_INPROC_SERVER+CLSCTX_LOCAL_SERVER)
#define CLSCTX_INPROC_HANDLER 2
#define CLSCTX_ALL (CLSCTX_INPROC_HANDLER+CLSCTX_INPROC_SERVER+CLSCTX_LOCAL_SERVER)
#define HIMETRIC_PER_INCH 2540
#define CFSTR_EMBEDSOURCE "Embed Source"
#define CFSTR_EMBEDDEDOBJECT "Embedded Object"
#define CFSTR_LINKSOURCE "Link Source"
#define CFSTR_CUSTOMLINKSOURCE "Custom Link Source"
#define CFSTR_OBJECTDESCRIPTOR "Object Descriptor"
#define CFSTR_LINKSRCDESCRIPTOR "Link Source Descriptor"
#define OLEUPDATE_ALWAYS 1
#define OLEUPDATE_ONCALL 3
#define OLELINKBIND_EVENIFCLASSDIFF 1
#define TKIND_ENUM 0
#define TKIND_RECORD (TKIND_ENUM + 1)
#define TKIND_MODULE (TKIND_RECORD + 1)
#define TKIND_INTERFACE (TKIND_MODULE + 1)
#define TKIND_DISPATCH (TKIND_INTERFACE + 1)
#define TKIND_COCLASS (TKIND_DISPATCH + 1)
#define TKIND_ALIAS (TKIND_COCLASS + 1)
#define TKIND_UNION (TKIND_ALIAS + 1)
#define TKIND_MAX (TKIND_UNION + 1)
#define DVASPECT_OPAQUE 16
#define DVASPECT_TRANSPARENT 32
#define DVASPECTINFOFLAG_CANOPTIMIZE 1
#define DISPATCH_METHOD 0x1
#define INVOKE_FUNC DISPATCH_METHOD
#define DISPID_UNKNOWN ( -1 )
#define MEMBERID_NIL DISPID_UNKNOWN
#define CC_FASTCALL 0
#define CC_CDECL 1
#define CC_MSCPASCAL (CC_CDECL + 1)
#define CC_PASCAL (CC_MSCPASCAL)
#define CC_MACPASCAL (CC_PASCAL + 1)
#define CC_STDCALL (CC_MACPASCAL + 1)
#define CC_FPFASTCALL (CC_STDCALL + 1)
#define CC_SYSCALL (CC_FPFASTCALL + 1)
#define CC_MPWCDECL (CC_SYSCALL + 1)
#define CC_MPWPASCAL (CC_MPWCDECL + 1)
#define CC_MAX (CC_MPWPASCAL + 1)
#define FUNC_VIRTUAL 0
#define FUNC_PUREVIRTUAL (FUNC_VIRTUAL + 1)
#define FUNC_NONVIRTUAL (FUNC_PUREVIRTUAL + 1)
#define FUNC_STATIC (FUNC_NONVIRTUAL + 1)
#define FUNC_DISPATCH (FUNC_STATIC + 1)
#define IMPLTYPEFLAG_FDEFAULT 0x1
#define IMPLTYPEFLAG_FSOURCE 0x2
#define IMPLTYPEFLAG_FRESTRICTED 0x4
#define IMPLTYPEFLAG_FDEFAULTVTABLE 0x800
#define VAR_PERINSTANCE 0
#define VAR_STATIC (VAR_PERINSTANCE+1)
#define VAR_CONST (VAR_STATIC+1)
#define VAR_DISPATCH (VAR_CONST+1)
#define OLEIVERB_PROPERTIES (-7)
#define STGM_DIRECT 0x00000000
#define STGM_TRANSACTED 0x00010000
#define STGM_SIMPLE 0x08000000
#define STGM_READ 0x00000000
#define STGM_WRITE 0x00000001
#define STGM_READWRITE 0x00000002
#define STGM_SHARE_DENY_NONE 0x00000040
#define STGM_SHARE_DENY_READ 0x00000030
#define STGM_SHARE_DENY_WRITE 0x00000020
#define STGM_SHARE_EXCLUSIVE 0x00000010
#define STGM_PRIORITY 0x00040000
#define STGM_DELETEONRELEASE 0x04000000
#define STGM_NOSCRATCH 0x00100000
#define STGM_CREATE 0x00001000
#define STGM_CONVERT 0x00020000
#define STGM_FAILIFTHERE 0x00000000
#define STGM_NOSNAPSHOT 0x00200000
#define ASYNC_MODE_COMPATIBILITY 0x00000001
#define ASYNC_MODE_DEFAULT 0x00000000
#define STGTY_REPEAT 0x00000100
#define STG_TOEND 0xFFFFFFFF
#define STG_LAYOUT_SEQUENTIAL 0x00000000
#define STG_LAYOUT_INTERLEAVED 0x00000001
#define STGFMT_STORAGE 0
#define STGFMT_NATIVE 1
#define STGFMT_FILE 3
#define STGFMT_ANY 4
#define STGFMT_DOCFILE 5
#define MKSYS_NONE 0
#define MKSYS_GENERICCOMPOSITE 1
#define MKSYS_FILEMONIKER 2
#define MKSYS_ANTIMONIKER 3
#define MKSYS_ITEMMONIKER 4
#define MKSYS_POINTERMONIKER 5
#define MKSYS_CLASSMONIKER 7
#define OLECLOSE_NOSAVE 1
#define OLECLOSE_PROMPTSAVE 2
#define OLECLOSE_SAVEIFDIRTY 0
#define OLEIVERB_DISCARDUNDOSTATE -6
#define OLEIVERB_HIDE -3
#define OLEIVERB_INPLACEACTIVATE -5
#define OLEIVERB_OPEN -2
#define OLEIVERB_PRIMARY 0
#define OLEIVERB_SHOW -1
#define OLEIVERB_UIACTIVATE -4
#define USERCLASSTYPE_APPNAME 3
#define USERCLASSTYPE_FULL 1
#define USERCLASSTYPE_SHORT 2
#define CONNECT_E_FIRST 0x80040200
#define CONNECT_E_ADVISELIMIT (CONNECT_E_FIRST+1)
#define CONNECT_E_CANNOTCONNECT (CONNECT_E_FIRST+2)
#define CONNECT_E_NOCONNECTION (CONNECT_E_FIRST+0)
#define CONNECT_E_OVERRIDDEN (CONNECT_E_FIRST+3)
#define STGTY_STORAGE 1
#define STGTY_STREAM 2
#define STGTY_LOCKBYTES 3
#define STGTY_PROPERTY 4
#define OLEUI_FALSE 0
#define OLEUI_SUCCESS 1
#define OLEUI_OK 1
#define OLEUI_CANCEL 2
#define OLEUI_ERR_STANDARDMIN 100
#define OLEUI_ERR_OLEMEMALLOC 100
#define OLEUI_ERR_STRUCTURENULL 101
#define OLEUI_ERR_STRUCTUREINVALID 102
#define OLEUI_ERR_CBSTRUCTINCORRECT 103
#define OLEUI_ERR_HWNDOWNERINVALID 104
#define OLEUI_ERR_LPSZCAPTIONINVALID 105
#define OLEUI_ERR_LPFNHOOKINVALID 106
#define OLEUI_ERR_HINSTANCEINVALID 107
#define OLEUI_ERR_LPSZTEMPLATEINVALID 108
#define OLEUI_ERR_HRESOURCEINVALID 109
#define OLEUI_ERR_FINDTEMPLATEFAILURE 110
#define OLEUI_ERR_LOADTEMPLATEFAILURE 111
#define OLEUI_ERR_DIALOGFAILURE 112
#define OLEUI_ERR_LOCALMEMALLOC 113
#define OLEUI_ERR_GLOBALMEMALLOC 114
#define OLEUI_ERR_LOADSTRING 115
#define OLEUI_ERR_STANDARDMAX 116
#define IOF_SHOWHELP 0x00000001L
#define IOF_SELECTCREATENEW 0x00000002L
#define IOF_SELECTCREATEFROMFILE 0x00000004L
#define IOF_CHECKLINK 0x00000008L
#define IOF_CHECKDISPLAYASICON 0x00000010L
#define IOF_CREATENEWOBJECT 0x00000020L
#define IOF_CREATEFILEOBJECT 0x00000040L
#define IOF_CREATELINKOBJECT 0x00000080L
#define IOF_DISABLELINK 0x00000100L
#define IOF_VERIFYSERVERSEXIST 0x00000200L
#define IOF_DISABLEDISPLAYASICON 0x00000400L
#define IOF_HIDECHANGEICON 0x00000800L
#define IOF_SHOWINSERTCONTROL 0x00001000L
#define IOF_SELECTCREATECONTROL 0x00002000L
#define OLEUI_IOERR_LPSZFILEINVALID (OLEUI_ERR_STANDARDMAX+0)
#define OLEUI_IOERR_LPSZLABELINVALID (OLEUI_ERR_STANDARDMAX+1)
#define OLEUI_IOERR_HICONINVALID (OLEUI_ERR_STANDARDMAX+2)
#define OLEUI_IOERR_LPFORMATETCINVALID (OLEUI_ERR_STANDARDMAX+3)
#define OLEUI_IOERR_PPVOBJINVALID (OLEUI_ERR_STANDARDMAX+4)
#define OLEUI_IOERR_LPIOLECLIENTSITEINVALID (OLEUI_ERR_STANDARDMAX+5)
#define OLEUI_IOERR_LPISTORAGEINVALID (OLEUI_ERR_STANDARDMAX+6)
#define OLEUI_IOERR_SCODEHASERROR (OLEUI_ERR_STANDARDMAX+7)
#define OLEUI_IOERR_LPCLSIDEXCLUDEINVALID (OLEUI_ERR_STANDARDMAX+8)
#define OLEUI_IOERR_CCHFILEINVALID (OLEUI_ERR_STANDARDMAX+9)
#define ODT_HEADER 100
#define ODT_TAB 101
#define ODT_LISTVIEW 102
#define LVM_FIRST 0x1000
#define TV_FIRST 0x1100
#define HDM_FIRST 0x1200
#define PGM_FIRST 0x1400
#define CCM_FIRST 0x2000
#define ECM_FIRST 0x1500
#define BCM_FIRST 0x1600
#define CBM_FIRST 0x1700
#define CCM_SETBKCOLOR (CCM_FIRST + 1)
#define CCM_SETCOLORSCHEME (CCM_FIRST + 2)
#define CCM_GETCOLORSCHEME (CCM_FIRST + 3)
#define CCM_GETDROPTARGET (CCM_FIRST + 4)
#define CCM_SETUNICODEFORMAT (CCM_FIRST + 5)
#define CCM_GETUNICODEFORMAT (CCM_FIRST + 6)
#define CCM_SETVERSION (CCM_FIRST + 0x7)
#define CCM_GETVERSION (CCM_FIRST + 0x8)
#define CCM_SETNOTIFYWINDOW (CCM_FIRST + 0x9)
#define CCM_SETWINDOWTHEME (CCM_FIRST + 0xb)
#define CCM_DPISCALE (CCM_FIRST + 0xc)
#define NM_FIRST (0U- 0U)
#define NM_LAST (0U- 99U)
#define NM_OUTOFMEMORY (NM_FIRST-1)
#define NM_CLICK (NM_FIRST-2)
#define NM_DBLCLK (NM_FIRST-3)
#define NM_RETURN (NM_FIRST-4)
#define NM_RCLICK (NM_FIRST-5)
#define NM_RDBLCLK (NM_FIRST-6)
#define NM_SETFOCUS (NM_FIRST-7)
#define NM_KILLFOCUS (NM_FIRST-8)
#define NM_CUSTOMDRAW (NM_FIRST-12)
#define NM_HOVER (NM_FIRST-13)
#define NM_NCHITTEST (NM_FIRST-14)
#define NM_KEYDOWN (NM_FIRST-15)
#define NM_RELEASEDCAPTURE (NM_FIRST-16)
#define NM_SETCURSOR (NM_FIRST-17)
#define NM_CHAR (NM_FIRST-18)
#define NM_TOOLTIPSCREATED (NM_FIRST-19)
#define NM_LDOWN (NM_FIRST-20)
#define NM_RDOWN (NM_FIRST-21)
#define NM_THEMECHANGED (NM_FIRST-22)
#define INFOTIPSIZE 1024
#define LVN_FIRST (0U-100U)
#define LVN_LAST (0U-199U)
#define HDN_FIRST (0U-300U)
#define HDN_LAST (0U-399U)
#define TVN_FIRST (0U-400U)
#define TVN_LAST (0U-499U)
#define TTN_FIRST (0U-520U)
#define TTN_LAST (0U-549U)
#define TCN_FIRST (0U-550U)
#define TCN_LAST (0U-580U)
#define CDN_FIRST (0U-601U)
#define CDN_LAST (0U-699U)
#define TBN_FIRST (0U-700U)
#define TBN_LAST (0U-720U)
#define UDN_FIRST (0U-721)
#define UDN_LAST (0U-740)
#define MSGF_COMMCTRL_BEGINDRAG 0x4200
#define MSGF_COMMCTRL_SIZEHEADER 0x4201
#define MSGF_COMMCTRL_DRAGSELECT 0x4202
#define MSGF_COMMCTRL_TOOLBARCUST 0x4203
#define CDRF_DODEFAULT 0x00000000
#define CDRF_NEWFONT 0x00000002
#define CDRF_SKIPDEFAULT 0x00000004
#define CDRF_NOTIFYPOSTPAINT 0x00000010
#define CDRF_NOTIFYITEMDRAW 0x00000020
#define CDRF_NOTIFYSUBITEMDRAW 0x00000020
#define CDRF_NOTIFYPOSTERASE 0x00000040
#define CDDS_PREPAINT 0x00000001
#define CDDS_POSTPAINT 0x00000002
#define CDDS_PREERASE 0x00000003
#define CDDS_POSTERASE 0x00000004
#define CDDS_ITEM 0x00010000
#define CDDS_ITEMPREPAINT 0x00010001
#define CDDS_ITEMPOSTPAINT 0x00010002
#define CDDS_ITEMPREERASE 0x00010003
#define CDDS_ITEMPOSTERASE 0x00010004
#define CDDS_SUBITEM 0x00020000
#define CDIS_SELECTED 0x0001
#define CDIS_GRAYED 0x0002
#define CDIS_DISABLED 0x0004
#define CDIS_CHECKED 0x0008
#define CDIS_FOCUS 0x0010
#define CDIS_DEFAULT 0x0020
#define CDIS_HOT 0x0040
#define CDIS_MARKED 0x0080
#define CDIS_INDETERMINATE 0x0100
#define CLR_NONE 0xFFFFFFFFL
#define CLR_DEFAULT 0xFF000000L
#define ILC_MASK 0x0001
#define ILC_COLOR 0x0000
#define ILC_COLORDDB 0x00FE
#define ILC_COLOR4 0x0004
#define ILC_COLOR8 0x0008
#define ILC_COLOR16 0x0010
#define ILC_COLOR24 0x0018
#define ILC_COLOR32 0x0020
#define ILC_PALETTE 0x0800
#define ILD_NORMAL 0x0000
#define ILD_TRANSPARENT 0x0001
#define ILD_MASK 0x0010
#define ILD_IMAGE 0x0020
#define ILD_BLEND25 0x0002
#define ILD_BLEND50 0x0004
#define ILD_OVERLAYMASK 0x0F00
#define ILD_SELECTED ILD_BLEND50
#define ILD_FOCUS ILD_BLEND25
#define ILD_BLEND ILD_BLEND50
#define CLR_HILIGHT CLR_DEFAULT
#define WC_HEADER "SysHeader32"
#define HDS_HORZ 0x00000000
#define HDS_BUTTONS 0x00000002
#define HDS_HOTTRACK 0x00000004
#define HDS_HIDDEN 0x00000008
#define HDS_DRAGDROP 0x00000040
#define HDS_FULLDRAG 0x00000080
#define HDS_FILTERBAR 0x00000100
#define HDS_FLAT 0x00000200
#define HDI_WIDTH 0x0001
#define HDI_HEIGHT HDI_WIDTH
#define HDI_TEXT 0x0002
#define HDI_FORMAT 0x0004
#define HDI_LPARAM 0x0008
#define HDI_BITMAP 0x0010
#define HDI_IMAGE 0x0020
#define HDI_DI_SETITEM 0x0040
#define HDI_ORDER 0x0080
#define HDI_FILTER 0x0100
#define HDF_LEFT 0
#define HDF_RIGHT 1
#define HDF_CENTER 2
#define HDF_JUSTIFYMASK 0x0003
#define HDF_RTLREADING 4
#define HDF_OWNERDRAW 0x8000
#define HDF_STRING 0x4000
#define HDF_BITMAP 0x2000
#define HDF_BITMAP_ON_RIGHT 0x1000
#define HDF_IMAGE 0x0800
#define HDF_SORTUP 0x0400
#define HDF_SORTDOWN 0x0200
#define HDM_GETITEMCOUNT (HDM_FIRST + 0)
#define HDM_INSERTITEMA (HDM_FIRST + 1)
#define HDM_INSERTITEMW (HDM_FIRST + 10)
#define HDM_INSERTITEM HDM_INSERTITEMA
#define HDM_DELETEITEM (HDM_FIRST + 2)
#define HDM_GETITEMA (HDM_FIRST + 3)
#define HDM_SETITEMA (HDM_FIRST + 4)
#define HDM_LAYOUT (HDM_FIRST + 5)
#define HDM_HITTEST (HDM_FIRST + 6)
#define HDM_GETITEMRECT (HDM_FIRST + 7)
#define HDM_SETIMAGELIST (HDM_FIRST + 8)
#define HDM_GETIMAGELIST (HDM_FIRST + 9)
#define HDM_GETITEMW (HDM_FIRST + 11)
#define HDM_SETITEMW (HDM_FIRST + 12)
#define HDM_ORDERTOINDEX (HDM_FIRST + 15)
#define HDM_CREATEDRAGIMAGE (HDM_FIRST + 16)
#define HDM_GETORDERARRAY (HDM_FIRST + 17)
#define HDM_SETORDERARRAY (HDM_FIRST + 18)
#define HDM_SETHOTDIVIDER (HDM_FIRST + 19)
#define HDM_GETITEM HDM_GETITEMA
#define HDM_SETITEM HDM_SETITEMA
#define HHT_NOWHERE 0x0001
#define HHT_ONHEADER 0x0002
#define HHT_ONDIVIDER 0x0004
#define HHT_ONDIVOPEN 0x0008
#define HHT_ONFILTER 0x0010
#define HHT_ONFILTERBUTTON 0x0020
#define HHT_ABOVE 0x0100
#define HHT_BELOW 0x0200
#define HHT_TORIGHT 0x0400
#define HHT_TOLEFT 0x0800
#define HDN_ITEMCHANGINGA (HDN_FIRST-0)
#define HDN_ITEMCHANGINGW (HDN_FIRST-20)
#define HDN_ITEMCHANGEDA (HDN_FIRST-1)
#define HDN_ITEMCHANGEDW (HDN_FIRST-21)
#define HDN_ITEMCLICKA (HDN_FIRST-2)
#define HDN_ITEMCLICKW (HDN_FIRST-22)
#define HDN_ITEMDBLCLICKA (HDN_FIRST-3)
#define HDN_ITEMDBLCLICKW (HDN_FIRST-23)
#define HDN_DIVIDERDBLCLICKA (HDN_FIRST-5)
#define HDN_DIVIDERDBLCLICKW (HDN_FIRST-25)
#define HDN_BEGINTRACKA (HDN_FIRST-6)
#define HDN_BEGINTRACKW (HDN_FIRST-26)
#define HDN_ENDTRACKA (HDN_FIRST-7)
#define HDN_ENDTRACKW (HDN_FIRST-27)
#define HDN_TRACKA (HDN_FIRST-8)
#define HDN_TRACKW (HDN_FIRST-28)
#define HDN_GETDISPINFOA (HDN_FIRST-9)
#define HDN_GETDISPINFOW (HDN_FIRST-29)
#define HDN_BEGINDRAG (HDN_FIRST-10)
#define HDN_ENDDRAG (HDN_FIRST-11)
#define HDN_FILTERCHANGE (HDN_FIRST-12)
#define HDN_FILTERBTNCLICK (HDN_FIRST-13)
#define HDN_ITEMCHANGING HDN_ITEMCHANGINGA
#define HDN_ITEMCHANGED HDN_ITEMCHANGEDA
#define HDN_ITEMCLICK HDN_ITEMCLICKA
#define HDN_ITEMDBLCLICK HDN_ITEMDBLCLICKA
#define HDN_DIVIDERDBLCLICK HDN_DIVIDERDBLCLICKA
#define HDN_BEGINTRACK HDN_BEGINTRACKA
#define HDN_ENDTRACK HDN_ENDTRACKA
#define HDN_TRACK HDN_TRACKA
#define TOOLBARCLASSNAME "ToolbarWindow32"
#define CMB_MASKED 0x02
#define TBSTATE_CHECKED 0x01
#define TBSTATE_PRESSED 0x02
#define TBSTATE_ENABLED 0x04
#define TBSTATE_HIDDEN 0x08
#define TBSTATE_INDETERMINATE 0x10
#define TBSTATE_WRAP 0x20
#define TBSTYLE_BUTTON 0x00
#define TBSTYLE_SEP 0x01
#define TBSTYLE_CHECK 0x02
#define TBSTYLE_GROUP 0x04
#define TBSTYLE_CHECKGROUP 0x06
#define TBSTYLE_TOOLTIPS 0x0100
#define TBSTYLE_WRAPABLE 0x0200
#define TBSTYLE_ALTDRAG 0x0400
#define WM_USER 0x0400
#define TB_ENABLEBUTTON (WM_USER + 1)
#define TB_CHECKBUTTON (WM_USER + 2)
#define TB_PRESSBUTTON (WM_USER + 3)
#define TB_HIDEBUTTON (WM_USER + 4)
#define TB_INDETERMINATE (WM_USER + 5)
#define TB_ISBUTTONENABLED (WM_USER + 9)
#define TB_ISBUTTONCHECKED (WM_USER + 10)
#define TB_ISBUTTONPRESSED (WM_USER + 11)
#define TB_ISBUTTONHIDDEN (WM_USER + 12)
#define TB_ISBUTTONINDETERMINATE (WM_USER + 13)
#define TB_SETSTATE (WM_USER + 17)
#define TB_GETSTATE (WM_USER + 18)
#define TB_ADDBITMAP (WM_USER + 19)
#define HINST_COMMCTRL PTR(_CAST, 0xFFFFFFFF)
#define IDB_STD_SMALL_COLOR 0
#define IDB_STD_LARGE_COLOR 1
#define IDB_VIEW_SMALL_COLOR 4
#define IDB_VIEW_LARGE_COLOR 5
#define IDB_HIST_SMALL_COLOR 8
#define IDB_HIST_LARGE_COLOR 9
#define STD_CUT 0
#define STD_COPY 1
#define STD_PASTE 2
#define STD_UNDO 3
#define STD_REDOW 4
#define STD_DELETE 5
#define STD_FILENEW 6
#define STD_FILEOPEN 7
#define STD_FILESAVE 8
#define STD_PRINTPRE 9
#define STD_PROPERTIES 10
#define STD_HELP 11
#define STD_FIND 12
#define STD_REPLACE 13
#define STD_PRINT 14
#define VIEW_LARGEICONS 0
#define VIEW_SMALLICONS 1
#define VIEW_LIST 2
#define VIEW_DETAILS 3
#define VIEW_SORTNAME 4
#define VIEW_SORTSIZE 5
#define VIEW_SORTDATE 6
#define VIEW_SORTTYPE 7
#define VIEW_PARENTFOLDER 8
#define VIEW_NETCONNECT 9
#define VIEW_NETDISCONNECT 10
#define VIEW_NEWFOLDER 11
#define VIEW_VIEWMENU 12
#define HIST_BACK 0
#define HIST_FORWARD 1
#define HIST_FAVORITES 2
#define HIST_ADDTOFAVORITES 3
#define HIST_VIEWTREE 4
#define TB_ADDBUTTONSA (WM_USER + 20)
#define TB_INSERTBUTTONA (WM_USER + 21)
#define TB_DELETEBUTTON (WM_USER + 22)
#define TB_GETBUTTON (WM_USER + 23)
#define TB_BUTTONCOUNT (WM_USER + 24)
#define TB_COMMANDTOINDEX (WM_USER + 25)
#define TB_SAVERESTOREA (WM_USER + 26)
#define TB_SAVERESTOREW (WM_USER + 76)
#define TB_CUSTOMIZE (WM_USER + 27)
#define TB_ADDSTRINGA (WM_USER + 28)
#define TB_ADDSTRINGW (WM_USER + 77)
#define TB_GETITEMRECT (WM_USER + 29)
#define TB_BUTTONSTRUCTSIZE (WM_USER + 30)
#define TB_SETBUTTONSIZE (WM_USER + 31)
#define TB_SETBITMAPSIZE (WM_USER + 32)
#define TB_AUTOSIZE (WM_USER + 33)
#define TB_GETTOOLTIPS (WM_USER + 35)
#define TB_SETTOOLTIPS (WM_USER + 36)
#define TB_SETPARENT (WM_USER + 37)
#define TB_SETROWS (WM_USER + 39)
#define TB_GETROWS (WM_USER + 40)
#define TB_GETBITMAPFLAGS (WM_USER + 41)
#define TB_SETCMDID (WM_USER + 42)
#define TB_CHANGEBITMAP (WM_USER + 43)
#define TB_GETBITMAP (WM_USER + 44)
#define TB_GETBUTTONTEXTA (WM_USER + 45)
#define TB_GETBUTTONTEXTW (WM_USER + 75)
#define TB_REPLACEBITMAP (WM_USER + 46)
#define TB_SETINDENT (WM_USER + 47)
#define TB_SETIMAGELIST (WM_USER + 48)
#define TB_GETIMAGELIST (WM_USER + 49)
#define TB_LOADIMAGES (WM_USER + 50)
#define TB_GETRECT (WM_USER + 51)
#define TB_SETHOTIMAGELIST (WM_USER + 52)
#define TB_GETHOTIMAGELIST (WM_USER + 53)
#define TB_SETDISABLEDIMAGELIST (WM_USER + 54)
#define TB_GETDISABLEDIMAGELIST (WM_USER + 55)
#define TB_SETSTYLE (WM_USER + 56)
#define TB_GETSTYLE (WM_USER + 57)
#define TB_GETBUTTONSIZE (WM_USER + 58)
#define TB_SETBUTTONWIDTH (WM_USER + 59)
#define TB_SETMAXTEXTROWS (WM_USER + 60)
#define TB_GETTEXTROWS (WM_USER + 61)
#define TB_GETBUTTONTEXT TB_GETBUTTONTEXTA
#define TB_SAVERESTORE TB_SAVERESTOREA
#define TB_ADDSTRING TB_ADDSTRINGA
#define TB_GETOBJECT (WM_USER + 62)
#define TB_GETHOTITEM (WM_USER + 71)
#define TB_SETHOTITEM (WM_USER + 72)
#define TB_SETANCHORHIGHLIGHT (WM_USER + 73)
#define TB_GETANCHORHIGHLIGHT (WM_USER + 74)
#define TB_MAPACCELERATORA (WM_USER + 78)
#define TBIMHT_AFTER 0x00000001
#define TBIMHT_BACKGROUND 0x00000002
#define TB_GETINSERTMARK (WM_USER + 79)
#define TB_SETINSERTMARK (WM_USER + 80)
#define TB_INSERTMARKHITTEST (WM_USER + 81)
#define TB_MOVEBUTTON (WM_USER + 82)
#define TB_GETMAXSIZE (WM_USER + 83)
#define TB_SETEXTENDEDSTYLE (WM_USER + 84)
#define TB_GETEXTENDEDSTYLE (WM_USER + 85)
#define TB_GETPADDING (WM_USER + 86)
#define TB_SETPADDING (WM_USER + 87)
#define TB_SETINSERTMARKCOLOR (WM_USER + 88)
#define TB_GETINSERTMARKCOLOR (WM_USER + 89)
#define TB_SETCOLORSCHEME CCM_SETCOLORSCHEME
#define TB_GETCOLORSCHEME CCM_GETCOLORSCHEME
#define TB_SETUNICODEFORMAT CCM_SETUNICODEFORMAT
#define TB_GETUNICODEFORMAT CCM_GETUNICODEFORMAT
#define TB_MAPACCELERATORW (WM_USER + 90)
#define TB_MAPACCELERATOR TB_MAPACCELERATORA
#define TBBF_LARGE 0x0001
#define TBIF_IMAGE 0x00000001
#define TBIF_TEXT 0x00000002
#define TBIF_STATE 0x00000004
#define TBIF_STYLE 0x00000008
#define TBIF_LPARAM 0x00000010
#define TBIF_COMMAND 0x00000020
#define TBIF_SIZE 0x00000040
#define TBIF_BYINDEX 0x80000000
#define TB_GETBUTTONINFOW (WM_USER + 63)
#define TB_SETBUTTONINFOW (WM_USER + 64)
#define TB_GETBUTTONINFOA (WM_USER + 65)
#define TB_SETBUTTONINFOA (WM_USER + 66)
#define TB_GETBUTTONINFO TB_GETBUTTONINFOA
#define TB_SETBUTTONINFO TB_SETBUTTONINFOA
#define TB_INSERTBUTTONW (WM_USER + 67)
#define TB_ADDBUTTONSW (WM_USER + 68)
#define TB_HITTEST (WM_USER + 69)
#define TB_INSERTBUTTON TB_INSERTBUTTONA
#define TB_ADDBUTTONS TB_ADDBUTTONSA
#define TB_SETDRAWTEXTFLAGS (WM_USER + 70)
#define TB_GETSTRINGW (WM_USER + 91)
#define TB_GETSTRINGA (WM_USER + 92)
#define TB_GETSTRING TB_GETSTRINGA
#define TBMF_PAD 0x00000001
#define TBMF_BARPAD 0x00000002
#define TBMF_BUTTONSPACING 0x00000004
#define TB_GETMETRICS (WM_USER + 101)
#define TB_SETMETRICS (WM_USER + 102)
#define TB_SETWINDOWTHEME CCM_SETWINDOWTHEME
#define TBN_GETBUTTONINFOA (TBN_FIRST-0)
#define TBN_GETBUTTONINFOW (TBN_FIRST-20)
#define TBN_BEGINDRAG (TBN_FIRST-1)
#define TBN_ENDDRAG (TBN_FIRST-2)
#define TBN_BEGINADJUST (TBN_FIRST-3)
#define TBN_ENDADJUST (TBN_FIRST-4)
#define TBN_RESET (TBN_FIRST-5)
#define TBN_QUERYINSERT (TBN_FIRST-6)
#define TBN_QUERYDELETE (TBN_FIRST-7)
#define TBN_TOOLBARCHANGE (TBN_FIRST-8)
#define TBN_CUSTHELP (TBN_FIRST-9)
#define TBN_DROPDOWN (TBN_FIRST - 10)
#define TBN_GETOBJECT (TBN_FIRST - 12)
#define TBN_GETBUTTONINFO TBN_GETBUTTONINFOA
#define TOOLTIPS_CLASS "tooltips_class32"
#define TTS_ALWAYSTIP 0x01
#define TTS_NOPREFIX 0x02
#define TTF_IDISHWND 0x01
#define TTF_CENTERTIP 0x02
#define TTF_RTLREADING 0x04
#define TTF_SUBCLASS 0x10
#define TTDT_AUTOMATIC 0
#define TTDT_RESHOW 1
#define TTDT_AUTOPOP 2
#define TTDT_INITIAL 3
#define TTM_ACTIVATE (WM_USER + 1)
#define TTM_SETDELAYTIME (WM_USER + 3)
#define TTM_ADDTOOL (WM_USER + 4)
#define TTM_ADDTOOLW (WM_USER + 50)
#define TTM_DELTOOL (WM_USER + 5)
#define TTM_DELTOOLW (WM_USER + 51)
#define TTM_NEWTOOLRECT (WM_USER + 6)
#define TTM_NEWTOOLRECTW (WM_USER + 52)
#define TTM_RELAYEVENT (WM_USER + 7)
#define TTM_GETTOOLINFO (WM_USER + 8)
#define TTM_GETTOOLINFOW (WM_USER + 53)
#define TTM_SETTOOLINFO (WM_USER + 9)
#define TTM_SETTOOLINFOW (WM_USER + 54)
#define TTM_HITTEST (WM_USER +10)
#define TTM_HITTESTW (WM_USER +55)
#define TTM_GETTEXT (WM_USER +11)
#define TTM_GETTEXTW (WM_USER +56)
#define TTM_UPDATETIPTEXT (WM_USER +12)
#define TTM_UPDATETIPTEXTW (WM_USER +57)
#define TTM_GETTOOLCOUNT (WM_USER +13)
#define TTM_ENUMTOOLS (WM_USER +14)
#define TTM_ENUMTOOLSW (WM_USER +58)
#define TTM_GETCURRENTTOOL (WM_USER + 15)
#define TTM_GETCURRENTTOOLW (WM_USER + 59)
#define TTM_winDOWFROMPOINT (WM_USER + 16)
#define TTN_NEEDTEXT (TTN_FIRST - 0)
#define TTN_NEEDTEXTW (TTN_FIRST - 10)
#define TTN_SHOW (TTN_FIRST - 1)
#define TTN_POP (TTN_FIRST - 2)
#define SBARS_SIZEGRIP 0x0100
#define STATUSCLASSNAME "msctls_statusbar32"
#define SB_SETTEXT (WM_USER+1)
#define SB_SETTEXTW (WM_USER+11)
#define SB_GETTEXT (WM_USER+2)
#define SB_GETTEXTW (WM_USER+13)
#define SB_GETTEXTLENGTH (WM_USER+3)
#define SB_GETTEXTLENGTHW (WM_USER+12)
#define SB_SETPARTS (WM_USER+4)
#define SB_GETPARTS (WM_USER+6)
#define SB_GETBORDERS (WM_USER+7)
#define SB_SETMINHEIGHT (WM_USER+8)
#define SB_SIMPLE (WM_USER+9)
#define SB_GETRECT (WM_USER+10)
#define SBT_OWNERDRAW 0x1000
#define SBT_NOBORDERS 0x0100
#define SBT_POPOUT 0x0200
#define SBT_RTLREADING 0x0400
#define SC_SIZE 0xF000
#define MINSYSCOMMAND SC_SIZE
#define TRACKBAR_CLASS "msctls_trackbar32"
#define TBS_AUTOTICKS 0x0001
#define TBS_VERT 0x0002
#define TBS_HORZ 0x0000
#define TBS_TOP 0x0004
#define TBS_BOTTOM 0x0000
#define TBS_LEFT 0x0004
#define TBS_RIGHT 0x0000
#define TBS_BOTH 0x0008
#define TBS_NOTICKS 0x0010
#define TBS_ENABLESELRANGE 0x0020
#define TBS_FIXEDLENGTH 0x0040
#define TBS_NOTHUMB 0x0080
#define TBS_TOOLTIPS 0x0100
#define TBM_GETPOS (WM_USER)
#define TBM_GETRANGEMIN (WM_USER+1)
#define TBM_GETRANGEMAX (WM_USER+2)
#define TBM_GETTIC (WM_USER+3)
#define TBM_SETTIC (WM_USER+4)
#define TBM_SETPOS (WM_USER+5)
#define TBM_SETRANGE (WM_USER+6)
#define TBM_SETRANGEMIN (WM_USER+7)
#define TBM_SETRANGEMAX (WM_USER+8)
#define TBM_CLEARTICS (WM_USER+9)
#define TBM_SETSEL (WM_USER+10)
#define TBM_SETSELSTART (WM_USER+11)
#define TBM_SETSELEND (WM_USER+12)
#define TBM_GETPTICS (WM_USER+14)
#define TBM_GETTICPOS (WM_USER+15)
#define TBM_GETNUMTICS (WM_USER+16)
#define TBM_GETSELSTART (WM_USER+17)
#define TBM_GETSELEND (WM_USER+18)
#define TBM_CLEARSEL (WM_USER+19)
#define TBM_SETTICFREQ (WM_USER+20)
#define TBM_SETPAGESIZE (WM_USER+21)
#define TBM_GETPAGESIZE (WM_USER+22)
#define TBM_SETLINESIZE (WM_USER+23)
#define TBM_GETLINESIZE (WM_USER+24)
#define TBM_GETTHUMBRECT (WM_USER+25)
#define TBM_GETCHANNELRECT (WM_USER+26)
#define TBM_SETTHUMBLENGTH (WM_USER+27)
#define TBM_GETTHUMBLENGTH (WM_USER+28)
#define TB_LINEUP 0
#define TB_LINEDOWN 1
#define TB_PAGEUP 2
#define TB_PAGEDOWN 3
#define TB_THUMBPOSITION 4
#define TB_THUMBTRACK 5
#define TB_TOP 6
#define TB_BOTTOM 7
#define TB_ENDTRACK 8
#define DL_BEGINDRAG (WM_USER+133)
#define DL_DRAGGING (WM_USER+134)
#define DL_DROPPED (WM_USER+135)
#define DL_CANCELDRAG (WM_USER+136)
#define DL_CURSORSET 0
#define DL_STOPCURSOR 1
#define DL_COPYCURSOR 2
#define DL_MOVECURSOR 3
#define DRAGLISTMSGSTRING "commctrl_DragListMsg"
#define UPDOWN_CLASS "msctls_updown32"
#define UD_MAXVAL 0x7fff
#define UD_MINVAL (-UD_MAXVAL)
#define UDS_WRAP 0x0001
#define UDS_SETBUDDYINT 0x0002
#define UDS_ALIGNRIGHT 0x0004
#define UDS_ALIGNLEFT 0x0008
#define UDS_AUTOBUDDY 0x0010
#define UDS_ARROWKEYS 0x0020
#define UDS_HORZ 0x0040
#define UDS_NOTHOUSANDS 0x0080
#define UDM_SETRANGE (WM_USER+101)
#define UDM_GETRANGE (WM_USER+102)
#define UDM_SETPOS (WM_USER+103)
#define UDM_GETPOS (WM_USER+104)
#define UDM_SETBUDDY (WM_USER+105)
#define UDM_GETBUDDY (WM_USER+106)
#define UDM_SETACCEL (WM_USER+107)
#define UDM_GETACCEL (WM_USER+108)
#define UDM_SETBASE (WM_USER+109)
#define UDM_GETBASE (WM_USER+110)
#define UDN_DELTAPOS (UDN_FIRST - 1)
#define PROGRESS_CLASS "msctls_progress32"
#define PBS_SMOOTH 0x01
#define PBS_VERTICAL 0x04
#define PBM_SETRANGE (WM_USER+1)
#define PBM_SETPOS (WM_USER+2)
#define PBM_DELTAPOS (WM_USER+3)
#define PBM_SETSTEP (WM_USER+4)
#define PBM_STEPIT (WM_USER+5)
#define PBM_SETRANGE32 (WM_USER+6)
#define PBM_GETRANGE (WM_USER+7)
#define PBM_GETPOS (WM_USER+8)
#define PBM_SETBARCOLOR (WM_USER+9)
#define PBM_SETBKCOLOR CCM_SETBKCOLOR
#define HOTKEYF_SHIFT 0x01
#define HOTKEYF_CONTROL 0x02
#define HOTKEYF_ALT 0x04
#define HOTKEYF_EXT 0x08
#define HKCOMB_NONE 0x0001
#define HKCOMB_S 0x0002
#define HKCOMB_C 0x0004
#define HKCOMB_A 0x0008
#define HKCOMB_SC 0x0010
#define HKCOMB_SA 0x0020
#define HKCOMB_CA 0x0040
#define HKCOMB_SCA 0x0080
#define HKM_SETHOTKEY (WM_USER+1)
#define HKM_GETHOTKEY (WM_USER+2)
#define HKM_SETRULES (WM_USER+3)
#define HOTKEY_CLASS "msctls_hotkey32"
#define CCS_TOP 0x00000001L
#define CCS_NOMOVEY 0x00000002L
#define CCS_BOTTOM 0x00000003L
#define CCS_NORESIZE 0x00000004L
#define CCS_NOPARENTALIGN 0x00000008L
#define CCS_ADJUSTABLE 0x00000020L
#define CCS_NODIVIDER 0x00000040L
#define WC_LISTVIEWA "SysListView32"
#define LVS_ICON 0x0000
#define LVS_REPORT 0x0001
#define LVS_SMALLICON 0x0002
#define LVS_LIST 0x0003
#define LVS_TYPEMASK 0x0003
#define LVS_SINGLESEL 0x0004
#define LVS_SHOWSELALWAYS 0x0008
#define LVS_SORTASCENDING 0x0010
#define LVS_SORTDESCENDING 0x0020
#define LVS_SHAREIMAGELISTS 0x0040
#define LVS_NOLABELWRAP 0x0080
#define LVS_AUTOARRANGE 0x0100
#define LVS_EDITLABELS 0x0200
#define LVS_OWNERDATA 0x1000
#define LVS_NOSCROLL 0x2000
#define LVS_TYPESTYLEMASK 0xfc00
#define LVS_ALIGNTOP 0x0000
#define LVS_ALIGNLEFT 0x0800
#define LVS_ALIGNMASK 0x0c00
#define LVS_OWNERDRAWFIXED 0x0400
#define LVS_NOCOLUMNHEADER 0x4000
#define LVS_NOSORTHEADER 0x8000
#define LVM_GETBKCOLOR (LVM_FIRST + 0)
#define LVM_SETBKCOLOR (LVM_FIRST + 1)
#define LVM_GETIMAGELIST (LVM_FIRST + 2)
#define LVSIL_NORMAL 0
#define LVSIL_SMALL 1
#define LVSIL_STATE 2
#define LVM_SETIMAGELIST (LVM_FIRST + 3)
#define LVM_GETITEMCOUNT (LVM_FIRST + 4)
#define LVIF_TEXT 0x0001
#define LVIF_IMAGE 0x0002
#define LVIF_PARAM 0x0004
#define LVIF_STATE 0x0008
#define LVIF_INDENT 0x0010
#define LVIF_NORECOMPUTE 0x0800
#define LVIS_FOCUSED 0x0001
#define LVIS_SELECTED 0x0002
#define LVIS_CUT 0x0004
#define LVIS_DROPHILITED 0x0008
#define LVIS_OVERLAYMASK 0x0F00
#define LVIS_STATEIMAGEMASK 0xF000
#define LPSTR_TEXTCALLBACK PSZ(_CAST, 0xFFFFFFFF)
#define I_IMAGECALLBACK (-1)
#define LVM_GETITEM (LVM_FIRST + 5)
#define LVM_SETITEM (LVM_FIRST + 6)
#define LVM_INSERTITEM (LVM_FIRST + 7)
#define LVM_DELETEITEM (LVM_FIRST + 8)
#define LVM_DELETEALLITEMS (LVM_FIRST + 9)
#define LVM_GETCALLBACKMASK (LVM_FIRST + 10)
#define LVM_SETCALLBACKMASK (LVM_FIRST + 11)
#define LVNI_ALL 0x0000
#define LVNI_FOCUSED 0x0001
#define LVNI_SELECTED 0x0002
#define LVNI_CUT 0x0004
#define LVNI_DROPHILITED 0x0008
#define LVNI_ABOVE 0x0100
#define LVNI_BELOW 0x0200
#define LVNI_TOLEFT 0x0400
#define LVNI_TORIGHT 0x0800
#define LVM_GETNEXTITEM (LVM_FIRST + 12)
#define LVFI_PARAM 0x0001
#define LVFI_STRING 0x0002
#define LVFI_PARTIAL 0x0008
#define LVFI_WRAP 0x0020
#define LVFI_NEARESTXY 0x0040
#define LVM_FINDITEM (LVM_FIRST + 13)
#define LVIR_BOUNDS 0
#define LVIR_ICON 1
#define LVIR_LABEL 2
#define LVIR_SELECTBOUNDS 3
#define LVM_GETITEMRECT (LVM_FIRST + 14)
#define LVM_SETITEMPOSITION (LVM_FIRST + 15)
#define LVM_GETITEMPOSITION (LVM_FIRST + 16)
#define LVM_GETSTRINGWIDTH (LVM_FIRST + 17)
#define LVHT_NOWHERE 0x0001
#define LVHT_ONITEMICON 0x0002
#define LVHT_ONITEMLABEL 0x0004
#define LVHT_ONITEMSTATEICON 0x0008
#define LVHT_ONITEM 0x000E
#define LVHT_ABOVE 0x0008
#define LVHT_BELOW 0x0010
#define LVHT_TORIGHT 0x0020
#define LVHT_TOLEFT 0x0040
#define LVM_HITTEST (LVM_FIRST + 18)
#define LVM_ENSUREVISIBLE (LVM_FIRST + 19)
#define LVM_SCROLL (LVM_FIRST + 20)
#define LVM_REDRAWITEMS (LVM_FIRST + 21)
#define LVA_DEFAULT 0x0000
#define LVA_ALIGNLEFT 0x0001
#define LVA_ALIGNTOP 0x0002
#define LVA_SNAPTOGRID 0x0005
#define LVM_ARRANGE (LVM_FIRST + 22)
#define LVM_EDITLABEL (LVM_FIRST + 23)
#define LVM_GETEDITCONTROL (LVM_FIRST + 24)
#define LVCF_FMT 0x0001
#define LVCF_WIDTH 0x0002
#define LVCF_TEXT 0x0004
#define LVCF_SUBITEM 0x0008
#define LVCFMT_LEFT 0x0000
#define LVCFMT_RIGHT 0x0001
#define LVCFMT_CENTER 0x0002
#define LVCFMT_JUSTIFYMASK 0x0003
#define LVM_GETCOLUMN (LVM_FIRST + 25)
#define LVM_SETCOLUMN (LVM_FIRST + 26)
#define LVM_INSERTCOLUMN (LVM_FIRST + 27)
#define LVM_DELETECOLUMN (LVM_FIRST + 28)
#define LVM_GETCOLUMNWIDTH (LVM_FIRST + 29)
#define LVSCW_AUTOSIZE -1
#define LVSCW_AUTOSIZE_USEHEADER -2
#define LVM_SETCOLUMNWIDTH (LVM_FIRST + 30)
#define LVM_CREATEDRAGIMAGE (LVM_FIRST + 33)
#define LVM_GETVIEWRECT (LVM_FIRST + 34)
#define LVM_GETTEXTCOLOR (LVM_FIRST + 35)
#define LVM_SETTEXTCOLOR (LVM_FIRST + 36)
#define LVM_GETTEXTBKCOLOR (LVM_FIRST + 37)
#define LVM_SETTEXTBKCOLOR (LVM_FIRST + 38)
#define LVM_GETTOPINDEX (LVM_FIRST + 39)
#define LVM_GETCOUNTPERPAGE (LVM_FIRST + 40)
#define LVM_GETORIGIN (LVM_FIRST + 41)
#define LVM_UPDATE (LVM_FIRST + 42)
#define LVM_SETITEMSTATE (LVM_FIRST + 43)
#define LVM_GETITEMSTATE (LVM_FIRST + 44)
#define LVM_GETITEMTEXT (LVM_FIRST + 45)
#define LVM_SETITEMTEXT (LVM_FIRST + 46)
#define LVSICF_NOINVALIDATEALL 0x00000001
#define LVSICF_NOSCROLL 0x00000002
#define LVM_SETITEMCOUNT (LVM_FIRST + 47)
#define LVM_SORTITEMS (LVM_FIRST + 48)
#define LVM_SETITEMPOSITION32 (LVM_FIRST + 49)
#define LVM_GETSELECTEDCOUNT (LVM_FIRST + 50)
#define LVM_GETITEMSPACING (LVM_FIRST + 51)
#define LVM_GETISEARCHSTRINGW (LVM_FIRST + 117)
#define LVM_GETISEARCHSTRING (LVM_FIRST + 52)
#define LVCDI_ITEM 0x00000000
#define LVCDI_GROUP 0x00000001
#define LVCDRF_NOSELECT 0x00010000
#define LVCDRF_NOGROUPFRAME 0x00020000
#define LVN_ITEMCHANGING (LVN_FIRST-0)
#define LVN_ITEMCHANGED (LVN_FIRST-1)
#define LVN_INSERTITEM (LVN_FIRST-2)
#define LVN_DELETEITEM (LVN_FIRST-3)
#define LVN_DELETEALLITEMS (LVN_FIRST-4)
#define LVN_BEGINLABELEDIT (LVN_FIRST-5)
#define LVN_BEGINLABELEDITW (LVN_FIRST-75)
#define LVN_ENDLABELEDIT (LVN_FIRST-6)
#define LVN_ENDLABELEDITW (LVN_FIRST-76)
#define LVN_COLUMNCLICK (LVN_FIRST-8)
#define LVN_BEGINDRAG (LVN_FIRST-9)
#define LVN_BEGINRDRAG (LVN_FIRST-11)
#define LVN_ODCACHEHINT (LVN_FIRST-13)
#define LVN_ODFINDITEM (LVN_FIRST-52)
#define LVN_ITEMACTIVATE (LVN_FIRST-14)
#define LVN_ODSTATECHANGED (LVN_FIRST-15)
#define LVN_GETDISPINFO (LVN_FIRST-50)
#define LVN_GETDISPINFOW (LVN_FIRST-77)
#define LVN_SETDISPINFO (LVN_FIRST-51)
#define LVN_SETDISPINFOW (LVN_FIRST-78)
#define LVIF_DI_SETITEM 0x1000
#define LVN_KEYDOWN (LVN_FIRST-55)
#define TVS_HASBUTTONS 0x0001
#define TVS_HASLINES 0x0002
#define TVS_LINESATROOT 0x0004
#define TVS_EDITLABELS 0x0008
#define TVS_DISABLEDRAGDROP 0x0010
#define TVS_SHOWSELALWAYS 0x0020
#define TVIF_TEXT 0x0001
#define TVIF_IMAGE 0x0002
#define TVIF_PARAM 0x0004
#define TVIF_STATE 0x0008
#define TVIF_HANDLE 0x0010
#define TVIF_SELECTEDIMAGE 0x0020
#define TVIF_CHILDREN 0x0040
#define TVIS_FOCUSED 0x0001
#define TVIS_SELECTED 0x0002
#define TVIS_CUT 0x0004
#define TVIS_DROPHILITED 0x0008
#define TVIS_BOLD 0x0010
#define TVIS_EXPANDED 0x0020
#define TVIS_EXPANDEDONCE 0x0040
#define TVIS_OVERLAYMASK 0x0F00
#define TVIS_STATEIMAGEMASK 0xF000
#define TVIS_USERMASK 0xF000
#define I_CHILDRENCALLBACK (-1)
#define TVI_ROOT PTR(_CAST, 0xFFFF0000)
#define TVI_FIRST PTR(_CAST, 0xFFFF0001)
#define TVI_LAST PTR(_CAST, 0xFFFF0002)
#define TVI_SORT PTR(_CAST, 0xFFFF0003)
#define TVM_INSERTITEM (TV_FIRST + 0)
#define TVM_DELETEITEM (TV_FIRST + 1)
#define TVM_EXPAND (TV_FIRST + 2)
#define TVE_COLLAPSE 0x0001
#define TVE_EXPAND 0x0002
#define TVE_TOGGLE 0x0003
#define TVE_COLLAPSERESET 0x8000
#define TVM_GETITEMRECT (TV_FIRST + 4)
#define TVM_GETCOUNT (TV_FIRST + 5)
#define TVM_GETINDENT (TV_FIRST + 6)
#define TVM_SETINDENT (TV_FIRST + 7)
#define TVM_GETIMAGELIST (TV_FIRST + 8)
#define TVSIL_NORMAL 0
#define TVSIL_STATE 2
#define TVM_SETIMAGELIST (TV_FIRST + 9)
#define TVM_GETNEXTITEM (TV_FIRST + 10)
#define TVGN_ROOT 0x0000
#define TVGN_NEXT 0x0001
#define TVGN_PREVIOUS 0x0002
#define TVGN_PARENT 0x0003
#define TVGN_CHILD 0x0004
#define TVGN_FIRSTVISIBLE 0x0005
#define TVGN_NEXTVISIBLE 0x0006
#define TVGN_PREVIOUSVISIBLE 0x0007
#define TVGN_DROPHILITE 0x0008
#define TVGN_CARET 0x0009
#define TVM_SELECTITEM (TV_FIRST + 11)
#define TVM_GETITEM (TV_FIRST + 12)
#define TVM_SETITEM (TV_FIRST + 13)
#define TVM_EDITLABEL (TV_FIRST + 14)
#define TVM_GETEDITCONTROL (TV_FIRST + 15)
#define TVM_GETVISIBLECOUNT (TV_FIRST + 16)
#define TVM_HITTEST (TV_FIRST + 17)
#define TVHT_NOWHERE 0x0001
#define TVHT_ONITEMICON 0x0002
#define TVHT_ONITEMLABEL 0x0004
#define TVHT_ONITEM 0x0046
#define TVHT_ONITEMINDENT 0x0008
#define TVHT_ONITEMBUTTON 0x0010
#define TVHT_ONITEMRIGHT 0x0020
#define TVHT_ONITEMSTATEICON 0x0040
#define TVHT_ABOVE 0x0100
#define TVHT_BELOW 0x0200
#define TVHT_TORIGHT 0x0400
#define TVHT_TOLEFT 0x0800
#define TVM_CREATEDRAGIMAGE (TV_FIRST + 18)
#define TVM_SORTCHILDREN (TV_FIRST + 19)
#define TVM_ENSUREVISIBLE (TV_FIRST + 20)
#define TVM_SORTCHILDRENCB (TV_FIRST + 21)
#define TVM_ENDEDITLABELNOW (TV_FIRST + 22)
#define TVM_GETISEARCHSTRING (TV_FIRST + 23)
#define TVN_SELCHANGINGA (TVN_FIRST-1)
#define TVN_SELCHANGINGW (TVN_FIRST-50)
#define TVN_SELCHANGEDA (TVN_FIRST-2)
#define TVN_SELCHANGEDW (TVN_FIRST-51)
#define TVC_UNKNOWN 0x0000
#define TVC_BYMOUSE 0x0001
#define TVC_BYKEYBOARD 0x0002
#define TVN_GETDISPINFOA (TVN_FIRST-3)
#define TVN_GETDISPINFOW (TVN_FIRST-52)
#define TVN_SETDISPINFOA (TVN_FIRST-4)
#define TVN_SETDISPINFOW (TVN_FIRST-53)
#define TVIF_DI_SETITEM 0x1000
#define TVN_ITEMEXPANDING (TVN_FIRST-5)
#define TVN_ITEMEXPANDED (TVN_FIRST-6)
#define TVN_BEGINDRAG (TVN_FIRST-7)
#define TVN_BEGINRDRAG (TVN_FIRST-8)
#define TVN_DELETEITEM (TVN_FIRST-9)
#define TVN_BEGINLABELEDIT (TVN_FIRST-10)
#define TVN_ENDLABELEDIT (TVN_FIRST-11)
#define TVN_KEYDOWN (TVN_FIRST-12)
#define WC_TABCONTROL "SysTabControl32"
#define TCS_SCROLLOPPOSITE 0x0001
#define TCS_BOTTOM 0x0002
#define TCS_RIGHT 0x0002
#define TCS_MULTISELECT 0x0004
#define TCS_FORCEICONLEFT 0x0010
#define TCS_FORCELABELLEFT 0x0020
#define TCS_HOTTRACK 0x0040
#define TCS_VERTICAL 0x0080
#define TCS_TABS 0x0000
#define TCS_BUTTONS 0x0100
#define TCS_SINGLELINE 0x0000
#define TCS_MULTILINE 0x0200
#define TCS_RIGHTJUSTIFY 0x0000
#define TCS_FIXEDWIDTH 0x0400
#define TCS_RAGGEDRIGHT 0x0800
#define TCS_FOCUSONBUTTONDOWN 0x1000
#define TCS_OWNERDRAWFIXED 0x2000
#define TCS_TOOLTIPS 0x4000
#define TCS_FOCUSNEVER 0x8000
#define TCM_FIRST 0x1300
#define TCM_GETIMAGELIST (TCM_FIRST + 2)
#define TCM_SETIMAGELIST (TCM_FIRST + 3)
#define TCM_GETITEMCOUNT (TCM_FIRST + 4)
#define TCIF_TEXT 0x0001
#define TCIF_IMAGE 0x0002
#define TCIF_RTLREADING 0x0004
#define TCIF_PARAM 0x0008
#define TCM_GETITEM (TCM_FIRST + 5)
#define TCM_SETITEM (TCM_FIRST + 6)
#define TCM_INSERTITEM (TCM_FIRST + 7)
#define TCM_DELETEITEM (TCM_FIRST + 8)
#define TCM_DELETEALLITEMS (TCM_FIRST + 9)
#define TCM_GETITEMRECT (TCM_FIRST + 10)
#define TCM_GETCURSEL (TCM_FIRST + 11)
#define TCM_SETCURSEL (TCM_FIRST + 12)
#define TCHT_NOWHERE 0x0001
#define TCHT_ONITEMICON 0x0002
#define TCHT_ONITEMLABEL 0x0004
#define TCHT_ONITEM 0x0006
#define TCM_HITTEST (TCM_FIRST + 13)
#define TCM_SETITEMEXTRA (TCM_FIRST + 14)
#define TCM_ADJUSTRECT (TCM_FIRST + 40)
#define TCM_SETITEMSIZE (TCM_FIRST + 41)
#define TCM_REMOVEIMAGE (TCM_FIRST + 42)
#define TCM_SETPADDING (TCM_FIRST + 43)
#define TCM_GETROWCOUNT (TCM_FIRST + 44)
#define TCM_GETTOOLTIPS (TCM_FIRST + 45)
#define TCM_SETTOOLTIPS (TCM_FIRST + 46)
#define TCM_GETCURFOCUS (TCM_FIRST + 47)
#define TCM_SETCURFOCUS (TCM_FIRST + 48)
#define TCN_KEYDOWN (TCN_FIRST - 0)
#define TCN_SELCHANGE (TCN_FIRST - 1)
#define TCN_SELCHANGING (TCN_FIRST - 2)
#define ANIMATE_CLASS "SysAnimate32"
#define ACS_CENTER 0x0001
#define ACS_TRANSPARENT 0x0002
#define ACS_AUTOPLAY 0x0004
#define ACM_OPENW (WM_USER+103)
#define ACM_OPEN (WM_USER+100)
#define ACM_PLAY (WM_USER+101)
#define ACM_STOP (WM_USER+102)
#define ACN_START 1
#define ACN_STOP 2
#define ICC_LISTVIEW_CLASSES 0x00000001
#define ICC_TREEVIEW_CLASSES 0x00000002
#define ICC_BAR_CLASSES 0x00000004
#define ICC_TAB_CLASSES 0x00000008
#define ICC_UPDOWN_CLASS 0x00000010
#define ICC_PROGRESS_CLASS 0x00000020
#define ICC_HOTKEY_CLASS 0x00000040
#define ICC_ANIMATE_CLASS 0x00000080
#define ICC_win95_CLASSES 0x000000FF
#define ICC_DATE_CLASSES 0x00000100
#define ICC_USEREX_CLASSES 0x00000200
#define ICC_COOL_CLASSES 0x00000400
#define ICC_INTERNET_CLASSES 0x00000800
#define ICC_PAGESCROLLER_CLASS 0x00001000
#define ICC_NATIVEFNTCTL_CLASS 0x00002000
#define ICC_STANDARD_CLASSES 0x00004000
#define ICC_LINK_CLASS 0x00008000
#define TBSTYLE_FLAT 0x0800
#define TTM_SETMAXTIPWIDTH (WM_USER + 24)
#define TTM_GETMAXTIPWIDTH (WM_USER + 25)
#define MCN_FIRST (0U-750U)
#define MCN_LAST (0U-759U)
#define MCM_FIRST 0x1000
#define MCM_GETCURSEL (MCM_FIRST + 1)
#define MCM_SETCURSEL (MCM_FIRST + 2)
#define MCM_GETMAXSELCOUNT (MCM_FIRST + 3)
#define MCM_SETMAXSELCOUNT (MCM_FIRST + 4)
#define MCM_GETSELRANGE (MCM_FIRST + 5)
#define MCM_SETSELRANGE (MCM_FIRST + 6)
#define MCM_GETMONTHRANGE (MCM_FIRST + 7)
#define MCM_SETDAYSTATE (MCM_FIRST + 8)
#define MCM_GETMINREQRECT (MCM_FIRST + 9)
#define MCM_SETTODAY (MCM_FIRST + 12)
#define MCM_GETTODAY (MCM_FIRST + 13)
#define MCM_HITTEST (MCM_FIRST + 14)
#define MCHT_TITLE 0x00010000
#define MCHT_CALENDAR 0x00020000
#define MCHT_TODAYLINK 0x00030000
#define MCHT_NEXT 0x01000000
#define MCHT_PREV 0x02000000
#define MCHT_NOWHERE 0x00000000
#define MCHT_TITLEBK 0x00010000
#define MCHT_TITLEMONTH 0x00010001
#define MCHT_TITLEYEAR 0x00010002
#define MCHT_TITLEBTNNEXT 0x01010003
#define MCHT_TITLEBTNPREV 0x02010003
#define MCHT_CALENDARBK 0x00020000
#define MCHT_CALENDARDATE 0x00020001
#define MCHT_CALENDARDATENEXT 0x01020001
#define MCHT_CALENDARDATEPREV 0x02020001
#define MCHT_CALENDARDAY 0x00020002
#define MCHT_CALENDARWEEKNUM 0x00020003
#define MCM_SETCOLOR (MCM_FIRST + 10)
#define MCM_GETCOLOR (MCM_FIRST + 11)
#define MCSC_BACKGROUND 0
#define MCSC_TEXT 1
#define MCSC_TITLEBK 2
#define MCSC_TITLETEXT 3
#define MCSC_MONTHBK 4
#define MCSC_TRAILINGTEXT 5
#define MCM_SETFIRSTDAYOFWEEK (MCM_FIRST + 15)
#define MCM_GETFIRSTDAYOFWEEK (MCM_FIRST + 16)
#define MCM_GETRANGE (MCM_FIRST + 17)
#define MCM_SETRANGE (MCM_FIRST + 18)
#define MCM_GETMONTHDELTA (MCM_FIRST + 19)
#define MCM_SETMONTHDELTA (MCM_FIRST + 20)
#define MCN_SELCHANGE (MCN_FIRST + 1)
#define MCN_GETDAYSTATE (MCN_FIRST + 3)
#define MCN_SELECT (MCN_FIRST + 4)
#define MCS_DAYSTATE 0x0001
#define MCS_MULTISELECT 0x0002
#define MCS_WEEKNUMBERS 0x0004
#define MCS_NOTODAYCIRCLE 0x0008
#define MCS_NOTODAY 0x0010
#define GMR_VISIBLE 0
#define GMR_DAYSTATE 1
#define DTN_FIRST (0U-760U)
#define DTN_LAST (0U-799U)
#define DTM_FIRST 0x1000
#define DTM_GETSYSTEMTIME (DTM_FIRST + 1)
#define DTM_SETSYSTEMTIME (DTM_FIRST + 2)
#define DTM_GETRANGE (DTM_FIRST + 3)
#define DTM_SETRANGE (DTM_FIRST + 4)
#define DTM_SETFORMAT (DTM_FIRST + 5)
#define DTM_SETMCCOLOR (DTM_FIRST + 6)
#define DTM_GETMCCOLOR (DTM_FIRST + 7)
#define DTM_GETMONTHCAL (DTM_FIRST + 8)
#define DTM_SETMCFONT (DTM_FIRST + 9)
#define DTM_GETMCFONT (DTM_FIRST + 10)
#define DTS_UPDOWN 0x0001
#define DTS_SHOWNONE 0x0002
#define DTS_SHORTDATEFORMAT 0x0000
#define DTS_LONGDATEFORMAT 0x0004
#define DTS_TIMEFORMAT 0x0009
#define DTS_APPCANPARSE 0x0010
#define DTS_RIGHTALIGN 0x0020
#define DTN_DATETIMECHANGE (DTN_FIRST + 1)
#define DTN_USERSTRING (DTN_FIRST + 2)
#define DTN_WMKEYDOWN (DTN_FIRST + 3)
#define DTN_FORMAT (DTN_FIRST + 4)
#define DTN_FORMATQUERY (DTN_FIRST + 5)
#define DTN_DROPDOWN (DTN_FIRST + 6)
#define DTN_CLOSEUP (DTN_FIRST + 7)
#define GDTR_MIN 0x0001
#define GDTR_MAX 0x0002
#define GDT_ERROR -1
#define GDT_VALID 0
#define GDT_NONE 1
#define LVM_SETEXTENDEDLISTVIEWSTYLE (LVM_FIRST + 54)
#define LVM_GETEXTENDEDLISTVIEWSTYLE (LVM_FIRST + 55)
#define LVS_EX_GRIDLINES 0x00000001
#define LVS_EX_SUBITEMIMAGES 0x00000002
#define LVS_EX_CHECKBOXES 0x00000004
#define LVS_EX_TRACKSELECT 0x00000008
#define LVS_EX_HEADERDRAGDROP 0x00000010
#define LVS_EX_FULLROWSELECT 0x00000020
#define LVS_EX_ONECLICKACTIVATE 0x00000040
#define LVS_EX_TWOCLICKACTIVATE 0x00000080
#define LVM_GETSUBITEMRECT (LVM_FIRST + 56)
#define LVM_SUBITEMHITTEST (LVM_FIRST + 57)
#define LVM_SETCOLUMNORDERARRAY (LVM_FIRST + 58)
#define LVM_GETCOLUMNORDERARRAY (LVM_FIRST + 59)
#define LVM_SETHOTITEM (LVM_FIRST + 60)
#define LVM_GETHOTITEM (LVM_FIRST + 61)
#define LVM_SETHOTCURSOR (LVM_FIRST + 62)
#define LVM_GETHOTCURSOR (LVM_FIRST + 63)
#define LVM_APPROXIMATEVIEWRECT (LVM_FIRST + 64)
#define LVM_SETWORKAREA (LVM_FIRST + 65)
#define RBIM_IMAGELIST 0x00000001
#define RBS_TOOLTIPS 0x0100
#define RBS_VARHEIGHT 0x0200
#define RBS_BANDBORDERS 0x0400
#define RBS_FIXEDORDER 0x0800
#define RBS_REGISTERDROP 0x1000
#define RBS_AUTOSIZE 0x2000
#define RBS_VERTICALGRIPPER 0x4000
#define RBS_DBLCLKTOGGLE 0x8000
#define RBBS_BREAK 0x00000001
#define RBBS_FIXEDSIZE 0x00000002
#define RBBS_CHILDEDGE 0x00000004
#define RBBS_HIDDEN 0x00000008
#define RBBS_NOVERT 0x00000010
#define RBBS_FIXEDBMP 0x00000020
#define RBBS_VARIABLEHEIGHT 0x00000040
#define RBBS_GRIPPERALWAYS 0x00000080
#define RBBS_NOGRIPPER 0x00000100
#define RBBIM_STYLE 0x00000001
#define RBBIM_COLORS 0x00000002
#define RBBIM_TEXT 0x00000004
#define RBBIM_IMAGE 0x00000008
#define RBBIM_CHILD 0x00000010
#define RBBIM_CHILDSIZE 0x00000020
#define RBBIM_SIZE 0x00000040
#define RBBIM_BACKGROUND 0x00000080
#define RBBIM_ID 0x00000100
#define RBBIM_IDEALSIZE 0x00000200
#define RBBIM_LPARAM 0x00000400
#define RBBIM_HEADERSIZE 0x00000800
#define RB_INSERTBAND (WM_USER + 1)
#define RB_DELETEBAND (WM_USER + 2)
#define RB_GETBARINFO (WM_USER + 3)
#define RB_SETBARINFO (WM_USER + 4)
#define RB_GETBANDINFO98 (WM_USER + 5)
#define RB_SETBANDINFO (WM_USER + 6)
#define RB_SETPARENT (WM_USER + 7)
#define RB_GETBANDCOUNT (WM_USER + 12)
#define RB_GETROWCOUNT (WM_USER + 13)
#define RB_GETROWHEIGHT (WM_USER + 14)
#define RB_HITTEST (WM_USER + 8)
#define RB_GETRECT (WM_USER + 9)
#define RB_IDTOINDEX (WM_USER + 16)
#define RB_GETTOOLTIPS (WM_USER + 17)
#define RB_SETTOOLTIPS (WM_USER + 18)
#define RB_SETBKCOLOR (WM_USER + 19)
#define RB_GETBKCOLOR (WM_USER + 20)
#define RB_SETTEXTCOLOR (WM_USER + 21)
#define RB_GETTEXTCOLOR (WM_USER + 22)
#define RB_SIZETORECT (WM_USER + 23)
#define RB_BEGINDRAG (WM_USER + 24)
#define RB_ENDDRAG (WM_USER + 25)
#define RB_DRAGMOVE (WM_USER + 26)
#define RB_GETBARHEIGHT (WM_USER + 27)
#define RB_GETBANDINFOW (WM_USER + 28)
#define RB_GETBANDINFOA (WM_USER + 29)
#define RB_GETBANDINFO RB_GETBANDINFOA
#define RB_MINIMIZEBAND (WM_USER + 30)
#define RB_MAXIMIZEBAND (WM_USER + 31)
#define RB_GETDROPTARGET (CCM_GETDROPTARGET)
#define RB_GETBANDBORDERS (WM_USER + 34)
#define RB_SHOWBAND (WM_USER + 35)
#define RB_SETPALETTE (WM_USER + 37)
#define RB_GETPALETTE (WM_USER + 38)
#define RB_MOVEBAND (WM_USER + 39)
#define RB_SETUNICODEFORMAT CCM_SETUNICODEFORMAT
#define RB_GETUNICODEFORMAT CCM_GETUNICODEFORMAT
#define RB_GETBANDMARGINS (WM_USER + 40)
#define RB_SETWINDOWTHEME CCM_SETWINDOWTHEME
#define RB_PUSHCHEVRON (WM_USER + 43)
#define RBN_FIRST (0U-831U)
#define RBN_LAST (0U-859U)
#define RBN_HEIGHTCHANGE (RBN_FIRST - 0)
#define RBN_GETOBJECT (RBN_FIRST - 1)
#define RBN_LAYOUTCHANGED (RBN_FIRST - 2)
#define RBN_AUTOSIZE (RBN_FIRST - 3)
#define RBN_BEGINDRAG (RBN_FIRST - 4)
#define RBN_ENDDRAG (RBN_FIRST - 5)
#define RBN_DELETINGBAND (RBN_FIRST - 6)
#define RBN_DELETEDBAND (RBN_FIRST - 7)
#define RBN_CHILDSIZE (RBN_FIRST - 8)
#define RBN_CHEVRONPUSHED (RBN_FIRST - 10)
#define RBN_MINMAX (RBN_FIRST - 21)
#define RBN_AUTOBREAK (RBN_FIRST - 22)
#define IPM_CLEARADDRESS (WM_USER+100)
#define IPM_SETADDRESS (WM_USER+101)
#define IPM_GETADDRESS (WM_USER+102)
#define IPM_SETRANGE (WM_USER+103)
#define IPM_SETFOCUS (WM_USER+104)
#define IPM_ISBLANK (WM_USER+105)
#define IPN_FIRST (0U-860U)
#define IPN_LAST (0U-879U)
#define IPN_FIELDCHANGED (IPN_FIRST - 0)
#define CBEIF_TEXT 0x00000001
#define CBEIF_IMAGE 0x00000002
#define CBEIF_SELECTEDIMAGE 0x00000004
#define CBEIF_OVERLAY 0x00000008
#define CBEIF_INDENT 0x00000010
#define CBEIF_LPARAM 0x00000020
#define CBEIF_DI_SETITEM 0x10000000
#define CBEM_INSERTITEM (WM_USER + 1)
#define CBEM_SETIMAGELIST (WM_USER + 2)
#define CBEM_GETIMAGELIST (WM_USER + 3)
#define CBEM_GETITEM (WM_USER + 4)
#define CBEM_SETITEM (WM_USER + 5)
#define CB_DELETESTRING 0x0144
#define CBEM_DELETEITEM CB_DELETESTRING
#define CBEM_GETCOMBOCONTROL (WM_USER + 6)
#define CBEM_GETEDITCONTROL (WM_USER + 7)
#define CBEM_SETEXSTYLE (WM_USER + 8)
#define CBEM_SETEXTENDEDSTYLE (WM_USER + 14)
#define CBEM_GETEXSTYLE (WM_USER + 9)
#define CBEM_HASEDITCHANGED (WM_USER + 10)
#define CBEM_INSERTITEMW (WM_USER + 11)
#define CBEM_SETITEMW (WM_USER + 12)
#define CBEM_GETITEMW (WM_USER + 13)
#define CBES_EX_NOEDITIMAGE 0x00000001
#define CBES_EX_NOEDITIMAGEINDENT 0x00000002
#define CBES_EX_PATHWORDBREAKPROC 0x00000004
#define CBES_EX_NOSIZELIMIT 0x00000008
#define CBES_EX_CASESENSITIVE 0x00000010
#define CBEN_FIRST (0U-800U)
#define CBEN_LAST (0U-830U)
#define CBEN_GETDISPINFO (CBEN_FIRST - 0)
#define CBEN_INSERTITEM (CBEN_FIRST - 1)
#define CBEN_DELETEITEM (CBEN_FIRST - 2)
#define CBEN_BEGINEDIT (CBEN_FIRST - 4)
#define CBEN_ENDEDIT (CBEN_FIRST - 5)
#define CBEN_DRAGBEGIN (CBEN_FIRST - 8)
#define CBENF_KILLFOCUS 1
#define CBENF_RETURN 2
#define CBENF_ESCAPE 3
#define CBENF_DROPDOWN 4
#define CBEMAXSTRLEN 260
#define BTNS_BUTTON TBSTYLE_BUTTON
#define BTNS_SEP TBSTYLE_SEP
#define BTNS_CHECK TBSTYLE_CHECK
#define BTNS_GROUP TBSTYLE_GROUP
#define BTNS_CHECKGROUP TBSTYLE_CHECKGROUP
#define TBSTYLE_DROPDOWN 0x0008
#define BTNS_DROPDOWN TBSTYLE_DROPDOWN
#define TBSTYLE_AUTOSIZE 0x0010
#define BTNS_AUTOSIZE TBSTYLE_AUTOSIZE
#define TBSTYLE_NOPREFIX 0x0020
#define BTNS_NOPREFIX TBSTYLE_NOPREFIX
#define BTNS_SHOWTEXT 0x0040
#define BTNS_WHOLEDROPDOWN 0x0080
#define TBSTYLE_EX_MIXEDBUTTONS 0x00000008
#define TBSTYLE_EX_HIDECLIPPEDBUTTONS 0x00000010
#define RBBS_USECHEVRON 0x00000200
#define RBBS_HIDETITLE 0x00000400
#define WMN_FIRST (0U-1000U)
#define WMN_LAST (0U-1200U)
#define RBHT_CHEVRON 0x0008
#define TTS_NOANIMATE 0x10
#define TTS_NOFADE 0x20
#define TTS_BALLOON 0x40
#define TTM_TRACKACTIVATE (WM_USER + 17)
#define TTM_TRACKPOSITION (WM_USER + 18)
#define TTM_SETTIPBKCOLOR (WM_USER + 19)
#define TTM_SETTIPTEXTCOLOR (WM_USER + 20)
#define TTM_GETDELAYTIME (WM_USER + 21)
#define TTM_GETTIPBKCOLOR (WM_USER + 22)
#define TTM_GETTIPTEXTCOLOR (WM_USER + 23)
#define TTM_SETMARGIN (WM_USER + 26)
#define TTM_GETMARGIN (WM_USER + 27)
#define TTM_POP (WM_USER + 28)
#define TTM_UPDATE (WM_USER + 29)
#define TTM_GETBUBBLESIZE (WM_USER + 30)
#define TTM_ADJUSTRECT (WM_USER + 31)
#define TTM_SETTITLEA (WM_USER + 32)
#define TTM_SETTITLEW (WM_USER + 33)
#define SBARS_TOOLTIPS 0x0800
#define UDM_SETRANGE32 (WM_USER+111)
#define UDM_GETRANGE32 (WM_USER+112)
#define UDM_SETUNICODEFORMAT CCM_SETUNICODEFORMAT
#define UDM_GETUNICODEFORMAT CCM_GETUNICODEFORMAT
#define UDM_SETPOS32 (WM_USER+113)
#define UDM_GETPOS32 (WM_USER+114)
#define LVS_EX_LABELTIP 0x00004000
#define TCN_GETOBJECT (TCN_FIRST - 3)
#define TCN_FOCUSCHANGE (TCN_FIRST - 4)
#define TBSTYLE_LIST 0x1000
#define TBSTYLE_CUSTOMERASE 0x2000
#define TBSTYLE_REGISTERDROP 0x4000
#define TBSTYLE_TRANSPARENT 0x8000
#define TBSTYLE_EX_DRAWDDARROWS 0x00000001
#define TBSTATE_ELLIPSES 0x40
#define TBSTATE_MARKED 0x80
#define SBN_FIRST (0U-880U)
#define SBN_LAST (0U-899U)
#define PGN_FIRST (0U-900U)
#define PGN_LAST (0U-950U)
#define TB_MARKBUTTON (WM_USER + 6)
#define TB_ISBUTTONHIGHLIGHTED (WM_USER + 14)
#define MAX_LINKID_TEXT 48
#define L_MAX_URL_LENGTH 2083
#define INVALID_LINK_INDEX (-1)
#define LWS_TRANSPARENT 0x0001
#define LWS_IGNORERETURN 0x0002
#define LIF_ITEMINDEX 0x00000001
#define LIF_STATE 0x00000002
#define LIF_ITEMID 0x00000004
#define LIF_URL 0x00000008
#define LIS_FOCUSED 0x00000001
#define LIS_ENABLED 0x00000002
#define LIS_VISITED 0x00000004
#define LM_HITTEST (WM_USER+0x300)
#define LM_GETIDEALHEIGHT (WM_USER+0x301)
#define LM_SETITEM (WM_USER+0x302)
#define LM_GETITEM (WM_USER+0x303)
#define LVGA_FOOTER_CENTER 0x00000010
#define LVGA_FOOTER_LEFT 0x00000008
#define LVGA_FOOTER_RIGHT 0x00000020
#define LVGA_HEADER_CENTER 0x00000002
#define LVGA_HEADER_LEFT 0x00000001
#define LVGA_HEADER_RIGHT 0x00000004
#define LVGF_ALIGN 0x00000008
#define LVGF_FOOTER 0x00000002
#define LVGF_GROUPID 0x00000010
#define LVGF_HEADER 0x00000001
#define LVGF_NONE 0x00000000
#define LVGF_STATE 0x00000004
#define LVGS_COLLAPSED 0x00000001
#define LVGS_HIDDEN 0x00000002
#define LVGS_NORMAL 0x00000000
#define LVIF_COLUMNS 0x0200
#define LVIF_GROUPID 0x0100
#define LVM_ENABLEGROUPVIEW (LVM_FIRST + 157)
#define LVM_GETGROUPINFO (LVM_FIRST + 148)
#define LVM_HASGROUP (LVM_FIRST + 161)
#define LVM_INSERTGROUP (LVM_FIRST + 145)
#define LVM_MOVEGROUP (LVM_FIRST + 151)
#define LVM_MOVEITEMTOGROUP (LVM_FIRST + 154)
#define LVM_REMOVEGROUP (LVM_FIRST + 150)
#define LVM_REMOVEALLGROUPS (LVM_FIRST + 160)
#define LVM_SETVIEW (LVM_FIRST + 142)
#define LV_VIEW_TILE 0x0004
#define LVM_ISGROUPVIEWENABLED (LVM_FIRST + 175)
#define LVM_SETGROUPINFO (LVM_FIRST + 147)
#define LVGMF_BORDERCOLOR 0x00000002
#define LVGMF_BORDERSIZE 0x00000001
#define LVGMF_NONE 0x00000000
#define LVGMF_TEXTCOLOR 0x00000004
#define LVM_SETGROUPMETRICS (LVM_FIRST + 155)
#define LVM_GETGROUPMETRICS (LVM_FIRST + 156)
#define LVBKIF_FLAG_TILEOFFSET 0x00000100
#define LVBKIF_SOURCE_HBITMAP 0x00000001
#define LVBKIF_SOURCE_MASK 0x00000003
#define LVBKIF_SOURCE_NONE 0x00000000
#define LVBKIF_SOURCE_URL 0x00000002
#define LVBKIF_STYLE_MASK 0x00000010
#define LVBKIF_STYLE_NORMAL 0x00000000
#define LVBKIF_STYLE_TILE 0x00000010
#define LVBKIF_TYPE_WATERMARK 0x10000000
#define LVM_GETBKIMAGEA (LVM_FIRST + 69)
#define LVM_GETBKIMAGEW (LVM_FIRST + 139)
#define LVM_GETHEADER (LVM_FIRST + 31)
#define LVM_GETSELECTEDCOLUMN (LVM_FIRST + 174)
#define LVM_SETBKIMAGEA (LVM_FIRST + 68)
#define LVM_SETBKIMAGE LVM_SETBKIMAGEA
#define LVM_SETBKIMAGEW (LVM_FIRST + 138)
#define LVM_SETSELECTEDCOLUMN (LVM_FIRST + 140)
#define LVS_EX_BORDERSELECT 0x00008000
#define LVS_EX_DOUBLEBUFFER 0x00010000
#define LVS_EX_HIDELABELS 0x00020000
#define LVS_EX_SIMPLESELECT 0x00100000
#define LVS_EX_SINGLEROW 0x00040000
#define LVS_EX_SNAPTOGRID 0x00080000
#define LV_VIEW_ICON 0x0000
#define LV_VIEW_DETAILS 0x0001
#define LV_VIEW_SMALLICON 0x0002
#define LV_VIEW_LIST 0x0003
#define HICF_OTHER 0x00000000
#define HICF_MOUSE 0x00000001
#define HICF_ARROWKEYS 0x00000002
#define HICF_ACCELERATOR 0x00000004
#define HICF_DUPACCEL 0x00000008
#define HICF_ENTERING 0x00000010
#define HICF_LEAVING 0x00000020
#define HICF_RESELECT 0x00000040
#define TBN_HOTITEMCHANGE (TBN_FIRST - 13)
#define TBN_DRAGOUT (TBN_FIRST - 14)
#define TBN_DELETINGBUTTON (TBN_FIRST - 15)
#define TBN_GETDISPINFOA (TBN_FIRST - 16)
#define TBN_GETDISPINFOW (TBN_FIRST - 17)
#define TBN_GETINFOTIPA (TBN_FIRST - 18)
#define TBN_GETINFOTIPW (TBN_FIRST - 19)
#define TBN_GETDISPINFO TBN_GETDISPINFOA
#define TBN_GETINFOTIP TBN_GETINFOTIPA
#define TBNF_IMAGE 0x00000001
#define TBNF_TEXT 0x00000002
#define TBNF_DI_SETITEM 0x10000000
#define TBDDRET_DEFAULT 0
#define TBDDRET_NODEFAULT 1
#define TBDDRET_TREATPRESSED 2
#define REBARCLASSNAME "ReBarWindow32"
#define TTF_TRACK 0x0020
#define TTF_ABSOLUTE 0x0080
#define TTF_TRANSPARENT 0x0100
#define TTF_DI_SETITEM 0x8000
#define SB_ISSIMPLE (WM_USER+14)
#define SB_SETICON (WM_USER+15)
#define SB_SETTIPTEXTA (WM_USER+16)
#define SB_SETTIPTEXTW (WM_USER+17)
#define SB_GETTIPTEXTA (WM_USER+18)
#define SB_GETTIPTEXTW (WM_USER+19)
#define SB_GETICON (WM_USER+20)
#define SB_SETTIPTEXT SB_SETTIPTEXTA
#define SB_GETTIPTEXT SB_GETTIPTEXTA
#define SBT_TOOLTIPS 0x0800
#define SBN_SIMPLEMODECHANGE (SBN_FIRST - 0)
#define TBM_SETTOOLTIPS (WM_USER+29)
#define TBM_GETTOOLTIPS (WM_USER+30)
#define TBM_SETTIPSIDE (WM_USER+31)
#define TBTS_TOP 0
#define TBTS_LEFT 1
#define TBTS_BOTTOM 2
#define TBTS_RIGHT 3
#define TBCD_TICS 0x0001
#define TBCD_THUMB 0x0002
#define TBCD_CHANNEL 0x0003
#define UDS_HOTTRACK 0x0100
#define CCS_VERT 0x00000080L
#define CCS_LEFT 0x00000081L
#define CCS_RIGHT 0x00000083L
#define CCS_NOMOVEX 0x00000082L
#define TBM_GETBUDDY (WM_USER+33)
#define LVCF_IMAGE 0x0010
#define LVCF_ORDER 0x0020
#define LVCFMT_IMAGE 0x0800
#define LVCFMT_BITMAP_ON_RIGHT 0x1000
#define LVCFMT_COL_HAS_IMAGES 0x8000
#define LVM_SETICONSPACING (LVM_FIRST + 53)
#define LV_MAX_WORKAREAS 16
#define LVM_SETWORKAREAS (LVM_FIRST + 65)
#define LVM_GETWORKAREAS (LVM_FIRST + 70)
#define LVM_GETNUMBEROFWORKAREAS (LVM_FIRST + 73)
#define LVM_GETSELECTIONMARK (LVM_FIRST + 66)
#define LVM_SETSELECTIONMARK (LVM_FIRST + 67)
#define LVM_SETHOVERTIME (LVM_FIRST + 71)
#define LVM_GETHOVERTIME (LVM_FIRST + 72)
#define LVM_SETTOOLTIPS (LVM_FIRST + 74)
#define LVM_GETTOOLTIPS (LVM_FIRST + 78)
#define LVM_GETBKIMAGE LVM_GETBKIMAGEA
#define LVKF_ALT 0x0001
#define LVKF_CONTROL 0x0002
#define LVKF_SHIFT 0x0004
#define LVN_HOTTRACK (LVN_FIRST-21)
#define LVN_ODFINDITEMA (LVN_FIRST-52)
#define LVN_ODFINDITEMW (LVN_FIRST-79)
#define LVN_GETDISPINFOA (LVN_FIRST-50)
#define LVN_SETDISPINFOA (LVN_FIRST-51)
#define LVN_MARQUEEBEGIN (LVN_FIRST-56)
#define LVGIT_UNFOLDED 0x0001
#define LVN_GETINFOTIPA (LVN_FIRST-57)
#define LVN_GETINFOTIPW (LVN_FIRST-58)
#define LVN_GETINFOTIP LVN_GETINFOTIPA
#define TVS_RTLREADING 0x0040
#define TVS_NOTOOLTIPS 0x0080
#define TVS_CHECKBOXES 0x0100
#define TVS_TRACKSELECT 0x0200
#define TVS_SINGLEEXPAND 0x0400
#define TVS_INFOTIP 0x0800
#define TVS_FULLROWSELECT 0x1000
#define TVS_NOSCROLL 0x2000
#define TVS_NONEVENHEIGHT 0x4000
#define TVS_NOHSCROLL 0x8000
#define TVIF_INTEGRAL 0x0080
#define TVIS_EXPANDPARTIAL 0x0080
#define TVE_EXPANDPARTIAL 0x4000
#define TVGN_LASTVISIBLE 0x000A
#define TVM_SETTOOLTIPS (TV_FIRST + 24)
#define TVM_GETTOOLTIPS (TV_FIRST + 25)
#define TVM_SETINSERTMARK (TV_FIRST + 26)
#define TVM_SETITEMHEIGHT (TV_FIRST + 27)
#define TVM_GETITEMHEIGHT (TV_FIRST + 28)
#define TVM_SETBKCOLOR (TV_FIRST + 29)
#define TVM_SETTEXTCOLOR (TV_FIRST + 30)
#define TVM_GETBKCOLOR (TV_FIRST + 31)
#define TVM_GETTEXTCOLOR (TV_FIRST + 32)
#define TVM_SETSCROLLTIME (TV_FIRST + 33)
#define TVM_GETSCROLLTIME (TV_FIRST + 34)
#define TVM_SETINSERTMARKCOLOR (TV_FIRST + 37)
#define TVM_GETINSERTMARKCOLOR (TV_FIRST + 38)
#define TVM_SETLINECOLOR (TV_FIRST + 40)
#define TVN_SELCHANGED TVN_SELCHANGEDA
#define TVN_GETDISPINFO TVN_GETDISPINFOA
#define TVN_GETINFOTIPA (TVN_FIRST-13)
#define TVN_GETINFOTIPW (TVN_FIRST-14)
#define TVN_SINGLEEXPAND (TVN_FIRST-15)
#define TVN_GETINFOTIP TVN_GETINFOTIPA
#define TVN_SELCHANGING TVN_SELCHANGINGA
#define TCS_EX_FLATSEPARATORS 0x00000001
#define TCS_EX_REGISTERDROP 0x00000002
#define TCIF_STATE 0x0010
#define TCIS_BUTTONPRESSED 0x0001
#define TCIS_HIGHLIGHTED 0x0002
#define TCM_HIGHLIGHTITEM (TCM_FIRST + 51)
#define TCM_SETEXTENDEDSTYLE (TCM_FIRST + 52)
#define TCM_GETEXTENDEDSTYLE (TCM_FIRST + 53)
#define ACS_TIMER 0x0008
#define RB_INSERTBANDA (WM_USER + 1)
#define RB_INSERTBANDW (WM_USER + 10)
#define RB_SETBANDINFOW (WM_USER + 11)
#define ILD_ROP 0x0040
#define FSB_REGULAR_MODE 0
#define FSB_ENCARTA_MODE 1
#define FSB_FLAT_MODE 2
#define MAXPROPPAGES 100
#define PSP_DEFAULT 0x00000000
#define PSP_DLGINDIRECT 0x00000001
#define PSP_USEHICON 0x00000002
#define PSP_USEICONID 0x00000004
#define PSP_USETITLE 0x00000008
#define PSP_RTLREADING 0x00000010
#define PSP_HASHELP 0x00000020
#define PSP_USEREFPARENT 0x00000040
#define PSP_USECALLBACK 0x00000080
#define PSP_PREMATURE 0x00000400
#define PSP_HIDEHEADER 0x00000800
#define PSP_USEHEADERTITLE 0x00001000
#define PSP_USEHEADERSUBTITLE 0x00002000
#define PSPCB_RELEASE 1
#define PSPCB_CREATE 2
#define PSH_DEFAULT 0x00000000
#define PSH_PROPTITLE 0x00000001
#define PSH_USEHICON 0x00000002
#define PSH_USEICONID 0x00000004
#define PSH_PROPSHEETPAGE 0x00000008
#define PSH_WIZARDHASFINISH 0x00000010
#define PSH_WIZARD 0x00000020
#define PSH_USEPSTARTPAGE 0x00000040
#define PSH_NOAPPLYNOW 0x00000080
#define PSH_USECALLBACK 0x00000100
#define PSH_HASHELP 0x00000200
#define PSH_MODELESS 0x00000400
#define PSH_RTLREADING 0x00000800
#define PSH_WIZARDCONTEXTHELP 0x00001000
#define PSH_WIZARD97 0x00002000
#define PSH_WATERMARK 0x00008000
#define PSH_USEHBMWATERMARK 0x00010000
#define PSH_USEHPLWATERMARK 0x00020000
#define PSH_STRETCHWATERMARK 0x00040000
#define PSH_HEADER 0x00080000
#define PSH_USEHBMHEADER 0x00100000
#define PSH_USEPAGELANG 0x00200000
#define PSCB_INITIALIZED 1
#define PSCB_PRECREATE 2
#define PSN_FIRST (0U-200U)
#define PSN_LAST (0U-299U)
#define PSN_SETACTIVE (PSN_FIRST-0)
#define PSN_KILLACTIVE (PSN_FIRST-1)
#define PSN_VALIDATE (PSN_FIRST-1)
#define PSN_APPLY (PSN_FIRST-2)
#define PSN_RESET (PSN_FIRST-3)
#define PSN_CANCEL (PSN_FIRST-3)
#define PSN_HELP (PSN_FIRST-5)
#define PSN_WIZBACK (PSN_FIRST-6)
#define PSN_WIZNEXT (PSN_FIRST-7)
#define PSN_WIZFINISH (PSN_FIRST-8)
#define PSN_QUERYCANCEL (PSN_FIRST-9)
#define PSN_GETOBJECT (PSN_FIRST-10)
#define PSNRET_NOERROR 0
#define PSNRET_INVALID 1
#define PSNRET_INVALID_NOCHANGEPAGE 2
#define PSM_SETCURSEL (WM_USER + 101)
#define PSM_REMOVEPAGE (WM_USER + 102)
#define PSM_ADDPAGE (WM_USER + 103)
#define PSM_CHANGED (WM_USER + 104)
#define PSM_RESTARTWINDOWS (WM_USER + 105)
#define PSM_REBOOTSYSTEM (WM_USER + 106)
#define PSM_CANCELTOCLOSE (WM_USER + 107)
#define PSM_QUERYSIBLINGS (WM_USER + 108)
#define PSM_UNCHANGED (WM_USER + 109)
#define PSM_APPLY (WM_USER + 110)
#define PSM_SETTITLEA (WM_USER + 111)
#define PSM_SETTITLEW (WM_USER + 120)
#define PSM_SETTITLE PSM_SETTITLEA
#define PSM_SETWIZBUTTONS (WM_USER + 112)
#define PSWIZB_BACK 0x00000001
#define PSWIZB_NEXT 0x00000002
#define PSWIZB_FINISH 0x00000004
#define PSWIZB_DISABLEDFINISH 0x00000008
#define PSM_PRESSBUTTON (WM_USER + 113)
#define PSBTN_BACK 0
#define PSBTN_NEXT 1
#define PSBTN_FINISH 2
#define PSBTN_OK 3
#define PSBTN_APPLYNOW 4
#define PSBTN_CANCEL 5
#define PSBTN_HELP 6
#define PSBTN_MAX 6
#define PSM_SETCURSELID (WM_USER + 114)
#define PSM_SETFINISHTEXTA (WM_USER + 115)
#define PSM_SETFINISHTEXTW (WM_USER + 121)
#define PSM_SETFINISHTEXT PSM_SETFINISHTEXTA
#define PSM_GETTABCONTROL (WM_USER + 116)
#define PSM_ISDIALOGMESSAGE (WM_USER + 117)
#define PSM_GETCURRENTPAGEHWND (WM_USER + 118)
#define ID_PSRESTARTWINDOWS 0x2
#define ID_PSREBOOTSYSTEM 0x3
#define PROP_SM_CXDLG 212
#define PROP_SM_CYDLG 188
#define PROP_MED_CXDLG 227
#define PROP_MED_CYDLG 215
#define PROP_LG_CXDLG 252
#define PROP_LG_CYDLG 218
#define WIZ_CXDLG 276
#define WIZ_CYDLG 140
#define WIZ_CXBMP 80
#define WIZ_BODYX 92
#define WIZ_BODYCX 184
#define WSB_PROP_CYVSCROLL 0x00000001L
#define WSB_PROP_CXHSCROLL 0x00000002L
#define WSB_PROP_CYHSCROLL 0x00000004L
#define WSB_PROP_CXVSCROLL 0x00000008L
#define WSB_PROP_CXHTHUMB 0x00000010L
#define WSB_PROP_CYVTHUMB 0x00000020L
#define WSB_PROP_VBKGCOLOR 0x00000040L
#define WSB_PROP_HBKGCOLOR 0x00000080L
#define WSB_PROP_VSTYLE 0x00000100L
#define WSB_PROP_HSTYLE 0x00000200L
#define WSB_PROP_winSTYLE 0x00000400L
#define WSB_PROP_PALETTE 0x00000800L
#define WSB_PROP_MASK 0x00000FFFL
#define TME_HOVER 0x00000001
#define TME_LEAVE 0x00000002
#define TME_QUERY 0x40000000
#define TME_CANCEL 0x80000000
#define HOVER_DEFAULT 0xFFFFFFFF
#define LVS_EX_FLATSB 0x00000100
#define LVS_EX_REGIONAL 0x00000200
#define LVS_EX_INFOTIP 0x00000400
#define LVS_EX_UNDERLINEHOT 0x00000800
#define LVS_EX_UNDERLINECOLD 0x00001000
#define OPENFILENAME_SIZE_VERSION_400 76
#define OFN_READONLY 0x00000001
#define OFN_OVERWRITEPROMPT 0x00000002
#define OFN_HIDEREADONLY 0x00000004
#define OFN_NOCHANGEDIR 0x00000008
#define OFN_SHOWHELP 0x00000010
#define OFN_ENABLEHOOK 0x00000020
#define OFN_ENABLETEMPLATE 0x00000040
#define OFN_ENABLETEMPLATEHANDLE 0x00000080
#define OFN_NOVALIDATE 0x00000100
#define OFN_ALLOWMULTISELECT 0x00000200
#define OFN_EXTENSIONDIFFERENT 0x00000400
#define OFN_PATHMUSTEXIST 0x00000800
#define OFN_FILEMUSTEXIST 0x00001000
#define OFN_CREATEPROMPT 0x00002000
#define OFN_SHAREAWARE 0x00004000
#define OFN_NOREADONLYRETURN 0x00008000
#define OFN_NOTESTFILECREATE 0x00010000
#define OFN_NONETWORKBUTTON 0x00020000
#define OFN_NOLONGNAMES 0x00040000
#define OFN_EXPLORER 0x00080000
#define OFN_NODEREFERENCELINKS 0x00100000
#define OFN_LONGNAMES 0x00200000
#define OFN_ENABLEINCLUDENOTIFY 0x00400000
#define OFN_ENABLESIZING 0x00800000
#define OFN_DONTADDTORECENT 0x02000000
#define OFN_FORCESHOWHIDDEN 0x10000000
#define OFN_SHAREFALLTHROUGH 2
#define OFN_SHARENOWARN 1
#define OFN_SHAREWARN 0
#define OFN_EX_NOPLACESBAR 0x00000001
#define CDN_INITDONE (CDN_FIRST - 0x0000)
#define CDN_SELCHANGE (CDN_FIRST - 0x0001)
#define CDN_FOLDERCHANGE (CDN_FIRST - 0x0002)
#define CDN_SHAREVIOLATION (CDN_FIRST - 0x0003)
#define CDN_HELP (CDN_FIRST - 0x0004)
#define CDN_FILEOK (CDN_FIRST - 0x0005)
#define CDN_TYPECHANGE (CDN_FIRST - 0x0006)
#define CDN_INCLUDEITEM (CDN_FIRST - 0x0007)
#define CDM_FIRST WM_USER +100
#define CDM_LAST WM_USER +200
#define CDM_GETSPEC (CDM_FIRST + 0x0000)
#define CDM_GETFILEPATH (CDM_FIRST + 0x0001)
#define CDM_GETFOLDERPATH (CDM_FIRST + 0x0002)
#define CDM_GETFOLDERIDLIST (CDM_FIRST + 0x0003)
#define CDM_SETCONTROLTEXT (CDM_FIRST + 0x0004)
#define CDM_HIDECONTROL (CDM_FIRST + 0x0005)
#define CDM_SETDEFEXT (CDM_FIRST + 0x0006)
#define CC_RGBINIT 0x00000001
#define CC_FULLOPEN 0x00000002
#define CC_PREVENTFULLOPEN 0x00000004
#define CC_SHOWHELP 0x00000008
#define CC_ENABLEHOOK 0x00000010
#define CC_ENABLETEMPLATE 0x00000020
#define CC_ENABLETEMPLATEHANDLE 0x00000040
#define CC_SOLIDCOLOR 0x00000080
#define CC_ANYCOLOR 0x00000100
#define FR_DOWN 0x00000001
#define FR_WHOLEWORD 0x00000002
#define FR_MATCHCASE 0x00000004
#define FR_FINDNEXT 0x00000008
#define FR_REPLACE 0x00000010
#define FR_REPLACEALL 0x00000020
#define FR_DIALOGTERM 0x00000040
#define FR_SHOWHELP 0x00000080
#define FR_ENABLEHOOK 0x00000100
#define FR_ENABLETEMPLATE 0x00000200
#define FR_NOUPDOWN 0x00000400
#define FR_NOMATCHCASE 0x00000800
#define FR_NOWHOLEWORD 0x00001000
#define FR_ENABLETEMPLATEHANDLE 0x00002000
#define FR_HIDEUPDOWN 0x00004000
#define FR_HIDEMATCHCASE 0x00008000
#define FR_HIDEWHOLEWORD 0x00010000
#define FR_RAW 0x00020000
#define FR_MATCHDIAC 0x20000000
#define FR_MATCHKASHIDA 0x40000000
#define FR_MATCHALEFHAMZA 0x80000000
#define CF_SCREENFONTS 0x00000001
#define CF_PRINTERFONTS 0x00000002
#define CF_BOTH 0x00000003
#define CF_SHOWHELP 0x00000004L
#define CF_ENABLEHOOK 0x00000008L
#define CF_ENABLETEMPLATE 0x00000010L
#define CF_ENABLETEMPLATEHANDLE 0x00000020L
#define CF_INITTOLOGFONTSTRUCT 0x00000040L
#define CF_USESTYLE 0x00000080L
#define CF_EFFECTS 0x00000100L
#define CF_APPLY 0x00000200L
#define CF_ANSIONLY 0x00000400L
#define CF_SCRIPTSONLY CF_ANSIONLY
#define CF_NOVECTORFONTS 0x00000800L
#define CF_NOOEMFONTS CF_NOVECTORFONTS
#define CF_NOSIMULATIONS 0x00001000L
#define CF_LIMITSIZE 0x00002000L
#define CF_FIXEDPITCHONLY 0x00004000L
#define CF_WYSIWYG 0x00008000L
#define CF_FORCEFONTEXIST 0x00010000L
#define CF_SCALABLEONLY 0x00020000L
#define CF_TTONLY 0x00040000L
#define CF_NOFACESEL 0x00080000L
#define CF_NOSTYLESEL 0x00100000L
#define CF_NOSIZESEL 0x00200000L
#define CF_SELECTSCRIPT 0x00400000L
#define CF_NOSCRIPTSEL 0x00800000L
#define CF_NOVERTFONTS 0x01000000L
#define SIMULATED_FONTTYPE 0x8000
#define PRINTER_FONTTYPE 0x4000
#define SCREEN_FONTTYPE 0x2000
#define BOLD_FONTTYPE 0x0100
#define ITALIC_FONTTYPE 0x0200
#define REGULAR_FONTTYPE 0x0400
#define PS_OPENTYPE_FONTTYPE 0x10000
#define TT_OPENTYPE_FONTTYPE 0x20000
#define TYPE1_FONTTYPE 0x40000
#define WM_CHOOSEFONT_GETLOGFONT (WM_USER + 1)
#define WM_CHOOSEFONT_SETLOGFONT (WM_USER + 101)
#define WM_CHOOSEFONT_SETFLAGS (WM_USER + 102)
#define LBSELCHSTRING "commdlg_LBSelChangedNotify"
#define SHAREVISTRING "commdlg_ShareViolation"
#define FILEOKSTRING "commdlg_FileNameOK"
#define COLOROKSTRING "commdlg_ColorOK"
#define SETRGBSTRING "commdlg_SetRGBColor"
#define HELPMSGSTRING "commdlg_help"
#define FINDMSGSTRING "commdlg_FindReplace"
#define CD_LBSELNOITEMS -1
#define CD_LBSELCHANGE 0
#define CD_LBSELSUB 1
#define CD_LBSELADD 2
#define PD_ALLPAGES 0x00000000
#define PD_SELECTION 0x00000001
#define PD_PAGENUMS 0x00000002
#define PD_NOSELECTION 0x00000004
#define PD_NOPAGENUMS 0x00000008
#define PD_COLLATE 0x00000010
#define PD_PRINTTOFILE 0x00000020
#define PD_PRINTSETUP 0x00000040
#define PD_NOWARNING 0x00000080
#define PD_RETURNDC 0x00000100
#define PD_RETURNIC 0x00000200
#define PD_RETURNDEFAULT 0x00000400
#define PD_SHOWHELP 0x00000800
#define PD_ENABLEPRINTHOOK 0x00001000
#define PD_ENABLESETUPHOOK 0x00002000
#define PD_ENABLEPRINTTEMPLATE 0x00004000
#define PD_ENABLESETUPTEMPLATE 0x00008000
#define PD_ENABLEPRINTTEMPLATEHANDLE 0x00010000
#define PD_ENABLESETUPTEMPLATEHANDLE 0x00020000
#define PD_USEDEVMODECOPIES 0x00040000
#define PD_USEDEVMODECOPIESANDCOLLATE 0x00040000
#define PD_DISABLEPRINTTOFILE 0x00080000
#define PD_HIDEPRINTTOFILE 0x00100000
#define PD_NONETWORKBUTTON 0x00200000
#define PD_CURRENTPAGE 0x00400000
#define PD_NOCURRENTPAGE 0x00800000
#define PD_EXCLUSIONFLAGS 0x01000000
#define PD_USELARGETEMPLATE 0x10000000
#define DM_COLLATE 0x00008000L
#define DM_COPIES 0x00000100L
#define PD_EXCL_COPIESANDCOLLATE (DM_COPIES | DM_COLLATE)
#define DN_DEFAULTPRN 0x0001
#define WM_PSD_PAGESETUPDLG (WM_USER )
#define WM_PSD_FULLPAGERECT (WM_USER+1)
#define WM_PSD_MINMARGINRECT (WM_USER+2)
#define WM_PSD_MARGINRECT (WM_USER+3)
#define WM_PSD_GREEKTEXTRECT (WM_USER+4)
#define WM_PSD_ENVSTAMPRECT (WM_USER+5)
#define WM_PSD_YAFULLPAGERECT (WM_USER+6)
#define PSD_DEFAULTMINMARGINS 0x00000000
#define PSD_INWININIINTLMEASURE 0x00000000
#define PSD_MINMARGINS 0x00000001
#define PSD_MARGINS 0x00000002
#define PSD_INTHOUSANDTHSOFINCHES 0x00000004
#define PSD_INHUNDREDTHSOFMILLIMETERS 0x00000008
#define PSD_DISABLEMARGINS 0x00000010
#define PSD_DISABLEPRINTER 0x00000020
#define PSD_NOWARNING 0x00000080
#define PSD_DISABLEORIENTATION 0x00000100
#define PSD_RETURNDEFAULT 0x00000400
#define PSD_DISABLEPAPER 0x00000200
#define PSD_SHOWHELP 0x00000800
#define PSD_ENABLEPAGESETUPHOOK 0x00002000
#define PSD_ENABLEPAGESETUPTEMPLATE 0x00008000
#define PSD_ENABLEPAGESETUPTEMPLATEHANDLE 0x00020000
#define PSD_ENABLEPAGEPAINTHOOK 0x00040000
#define PSD_DISABLEPAGEPAINTING 0x00080000
#define PSD_NONETWORKBUTTON 0x00200000
#define _UPPER 0x1
#define _LOWER 0x2
#define _DIGIT 0x4
#define _SPACE 0x8
#define _PUNCT 0x10
#define _CONTROL 0x20
#define _BLANK 0x40
#define __HEX 0x80
#define _LEADBYTE 0x8000
#define _ALPHA 0x0103
#define WM_DDE_FIRST 0x03E0
#define WM_DDE_INITIATE (WM_DDE_FIRST)
#define WM_DDE_TERMINATE (WM_DDE_FIRST+1)
#define WM_DDE_ADVISE (WM_DDE_FIRST+2)
#define WM_DDE_UNADVISE (WM_DDE_FIRST+3)
#define WM_DDE_ACK (WM_DDE_FIRST+4)
#define WM_DDE_DATA (WM_DDE_FIRST+5)
#define WM_DDE_REQUEST (WM_DDE_FIRST+6)
#define WM_DDE_POKE (WM_DDE_FIRST+7)
#define WM_DDE_EXECUTE (WM_DDE_FIRST+8)
#define WM_DDE_LAST (WM_DDE_FIRST+8)
#define XST_NULL 0
#define XST_INCOMPLETE 1
#define XST_CONNECTED 2
#define XST_INIT1 3
#define XST_INIT2 4
#define XST_REQSENT 5
#define XST_DATARCVD 6
#define XST_POKESENT 7
#define XST_POKEACKRCVD 8
#define XST_EXECSENT 9
#define XST_EXECACKRCVD 10
#define XST_ADVSENT 11
#define XST_UNADVSENT 12
#define XST_ADVACKRCVD 13
#define XST_UNADVACKRCVD 14
#define XST_ADVDATASENT 15
#define XST_ADVDATAACKRCVD 16
#define CADV_LATEACK 0xFFFF
#define ST_CONNECTED 0x0001
#define ST_ADVISE 0x0002
#define ST_ISLOCAL 0x0004
#define ST_BLOCKED 0x0008
#define ST_CLIENT 0x0010
#define ST_TERMINATED 0x0020
#define ST_INLIST 0x0040
#define ST_BLOCKNEXT 0x0080
#define ST_ISSELF 0x0100
#define DDE_FACK 0x8000
#define DDE_FBUSY 0x4000
#define DDE_FDEFERUPD 0x4000
#define DDE_FACKREQ 0x8000
#define DDE_FRELEASE 0x2000
#define DDE_FREQUESTED 0x1000
#define DDE_FAPPSTATUS 0x00ff
#define DDE_FNOTPROCESSED 0x0000
#define DDE_FACKRESERVED 0x3F00
#define DDE_FADVRESERVED 0X3FFF
#define DDE_FDATRESERVED 0X4FFF
#define DDE_FPOKRESERVED 0xDFFF
#define MSGF_DDEMGR 0x8001
#define CP_WINANSI 1004
#define CP_WINUNICODE 1200
#define XTYPF_NOBLOCK 0x0002
#define XTYPF_NODATA 0x0004
#define XTYPF_ACKREQ 0x0008
#define XCLASS_MASK 0xFC00
#define XCLASS_BOOL 0x1000
#define XCLASS_DATA 0x2000
#define XCLASS_FLAGS 0x4000
#define XCLASS_NOTIFICATION 0x8000
#define XTYP_ERROR 0x8002
#define XTYP_ADVDATA 0x4010
#define XTYP_ADVREQ 0x2022
#define XTYP_ADVSTART 0x1030
#define XTYP_ADVSTOP 0x8040
#define XTYP_EXECUTE 0x4050
#define XTYP_CONNECT 0x1062
#define XTYP_CONNECT_CONFIRM 0x8072
#define XTYP_XACT_COMPLETE 0x8080
#define XTYP_POKE 0x4090
#define XTYP_REGISTER 0x80A2
#define XTYP_REQUEST 0x20B0
#define XTYP_DISCONNECT 0x80c2
#define XTYP_UNREGISTER 0x80d2
#define XTYP_WILDCONNECT 0x20e2
#define XTYP_MASK 0x00F0
#define XTYP_SHIFT 4
#define TIMEOUT_ASYNC 0xFFFFFFFF
#define QID_SYNC 0xFFFFFFFF
#define SZDDESYS_TOPIC "System"
#define SZDDESYS_ITEM_TOPICS "Topics"
#define SZDDESYS_ITEM_SYSITEMS "SysItems"
#define SZDDESYS_ITEM_RTNMSG "ReturnMessage"
#define SZDDESYS_ITEM_STATUS "Status"
#define SZDDESYS_ITEM_FORMATS "Formats"
#define SZDDESYS_ITEM_HELP "Help"
#define SZDDE_ITEM_ITEMLIST "TopicItemList"
#define CBR_BLOCK ptr(_cast, 0xffffffffL)
#define CBF_FAIL_SELFCONNECTIONS 0x00001000
#define CBF_FAIL_CONNECTIONS 0x00002000
#define CBF_FAIL_ADVISES 0x00004000
#define CBF_FAIL_EXECUTES 0x00008000
#define CBF_FAIL_POKES 0x00010000
#define CBF_FAIL_REQUESTS 0x00020000
#define CBF_FAIL_ALLSVRXACTIONS 0x0003f000
#define CBF_SKIP_CONNECT_CONFIRMS 0x00040000
#define CBF_SKIP_REGISTRATIONS 0x00080000
#define CBF_SKIP_UNREGISTRATIONS 0x00100000
#define CBF_SKIP_DISCONNECTS 0x00200000
#define CBF_SKIP_ALLNOTIFICATIONS 0x003c0000
#define APPCMD_CLIENTONLY 0x00000010L
#define APPCMD_FILTERINITS 0x00000020L
#define APPCMD_MASK 0x00000FF0L
#define APPCLASS_STANDARD 0x00000000L
#define APPCLASS_MASK 0x0000000FL
#define EC_ENABLEALL 0
#define EC_ENABLEONE ST_BLOCKNEXT
#define EC_DISABLE ST_BLOCKED
#define EC_QUERYWAITING 2
#define DNS_REGISTER 0x0001
#define DNS_UNREGISTER 0x0002
#define DNS_FILTERON 0x0004
#define DNS_FILTEROFF 0x0008
#define HDATA_APPOWNED 0x0001
#define DMLERR_NO_ERROR 0
#define DMLERR_FIRST 0x4000
#define DMLERR_ADVACKTIMEOUT 0x4000
#define DMLERR_BUSY 0x4001
#define DMLERR_DATAACKTIMEOUT 0x4002
#define DMLERR_DLL_NOT_INITIALIZED 0x4003
#define DMLERR_DLL_USAGE 0x4004
#define DMLERR_EXECACKTIMEOUT 0x4005
#define DMLERR_INVALIDPARAMETER 0x4006
#define DMLERR_LOW_MEMORY 0x4007
#define DMLERR_MEMORY_ERROR 0x4008
#define DMLERR_NOTPROCESSED 0x4009
#define DMLERR_NO_CONV_ESTABLISHED 0x400a
#define DMLERR_POKEACKTIMEOUT 0x400b
#define DMLERR_POSTMSG_FAILED 0x400c
#define DMLERR_REENTRANCY 0x400d
#define DMLERR_SERVER_DIED 0x400e
#define DMLERR_SYS_ERROR 0x400f
#define DMLERR_UNADVACKTIMEOUT 0x4010
#define DMLERR_UNFOUND_QUEUE_ID 0x4011
#define DMLERR_LAST 0x4011
#define MH_CREATE 1
#define MH_KEEP 2
#define MH_DELETE 3
#define MH_CLEANUP 4
#define MAX_MONITORS 4
#define APPCLASS_MONITOR 0x00000001L
#define XTYP_MONITOR 0x000080F2L
#define MF_HSZ_INFO 0x01000000
#define MF_SENDMSGS 0x02000000
#define MF_POSTMSGS 0x04000000
#define MF_CALLBACKS 0x08000000
#define MF_ERRORS 0x10000000
#define MF_LINKS 0x20000000
#define MF_CONV 0x40000000
#define MF_MASK 0xFF000000
#define ctlFirst 0x0400
#define ctlLast 0x04ff
#define psh1 0x0400
#define psh2 0x0401
#define psh3 0x0402
#define psh4 0x0403
#define psh5 0x0404
#define psh6 0x0405
#define psh7 0x0406
#define psh8 0x0407
#define psh9 0x0408
#define psh10 0x0409
#define psh11 0x040a
#define psh12 0x040b
#define psh13 0x040c
#define psh14 0x040d
#define psh15 0x040e
#define pshHelp psh15
#define psh16 0x040f
#define chx1 0x0410
#define chx2 0x0411
#define chx3 0x0412
#define chx4 0x0413
#define chx5 0x0414
#define chx6 0x0415
#define chx7 0x0416
#define chx8 0x0417
#define chx9 0x0418
#define chx10 0x0419
#define chx11 0x041a
#define chx12 0x041b
#define chx13 0x041c
#define chx14 0x041d
#define chx15 0x041e
#define chx16 0x041f
#define rad1 0x0420
#define rad2 0x0421
#define rad3 0x0422
#define rad4 0x0423
#define rad5 0x0424
#define rad6 0x0425
#define rad7 0x0426
#define rad8 0x0427
#define rad9 0x0428
#define rad10 0x0429
#define rad11 0x042a
#define rad12 0x042b
#define rad13 0x042c
#define rad14 0x042d
#define rad15 0x042e
#define rad16 0x042f
#define grp1 0x0430
#define grp2 0x0431
#define grp3 0x0432
#define grp4 0x0433
#define frm1 0x0434
#define frm2 0x0435
#define frm3 0x0436
#define frm4 0x0437
#define rct1 0x0438
#define rct2 0x0439
#define rct3 0x043a
#define rct4 0x043b
#define ico1 0x043c
#define ico2 0x043d
#define ico3 0x043e
#define ico4 0x043f
#define stc1 0x0440
#define stc2 0x0441
#define stc3 0x0442
#define stc4 0x0443
#define stc5 0x0444
#define stc6 0x0445
#define stc7 0x0446
#define stc8 0x0447
#define stc9 0x0448
#define stc10 0x0449
#define stc11 0x044a
#define stc12 0x044b
#define stc13 0x044c
#define stc14 0x044d
#define stc15 0x044e
#define stc16 0x044f
#define stc17 0x0450
#define stc18 0x0451
#define stc19 0x0452
#define stc20 0x0453
#define stc21 0x0454
#define stc22 0x0455
#define stc23 0x0456
#define stc24 0x0457
#define stc25 0x0458
#define stc26 0x0459
#define stc27 0x045a
#define stc28 0x045b
#define stc29 0x045c
#define stc30 0x045d
#define stc31 0x045e
#define stc32 0x045f
#define lst1 0x0460
#define lst2 0x0461
#define lst3 0x0462
#define lst4 0x0463
#define lst5 0x0464
#define lst6 0x0465
#define lst7 0x0466
#define lst8 0x0467
#define lst9 0x0468
#define lst10 0x0469
#define lst11 0x046a
#define lst12 0x046b
#define lst13 0x046c
#define lst14 0x046d
#define lst15 0x046e
#define lst16 0x046f
#define cmb1 0x0470
#define cmb2 0x0471
#define cmb3 0x0472
#define cmb4 0x0473
#define cmb5 0x0474
#define cmb6 0x0475
#define cmb7 0x0476
#define cmb8 0x0477
#define cmb9 0x0478
#define cmb10 0x0479
#define cmb11 0x047a
#define cmb12 0x047b
#define cmb13 0x047c
#define cmb14 0x047d
#define cmb15 0x047e
#define cmb16 0x047f
#define edt1 0x0480
#define edt2 0x0481
#define edt3 0x0482
#define edt4 0x0483
#define edt5 0x0484
#define edt6 0x0485
#define edt7 0x0486
#define edt8 0x0487
#define edt9 0x0488
#define edt10 0x0489
#define edt11 0x048a
#define edt12 0x048b
#define edt13 0x048c
#define edt14 0x048d
#define edt15 0x048e
#define edt16 0x048f
#define scr1 0x0490
#define scr2 0x0491
#define scr3 0x0492
#define scr4 0x0493
#define scr5 0x0494
#define scr6 0x0495
#define scr7 0x0496
#define scr8 0x0497
#define ctl1 0x04A0
#define FILEOPENORD 1536
#define MULTIFILEOPENORD 1537
#define PRINTDLGORD 1538
#define PRNSETUPDLGORD 1539
#define FINDDLGORD 1540
#define REPLACEDLGORD 1541
#define FONTDLGORD 1542
#define FORMATDLGORD31 1543
#define FORMATDLGORD30 1544
#define RUNDLGORD 1545
#define PAGESETUPDLGORD 1546
#define NEWFILEOPENORD 1547
#define PRINTDLGEXORD 1549
#define PAGESETUPDLGORDMOTIF 1550
#define COLORMGMTDLGORD 1551
#define NEWFILEOPENV2ORD 1552
#define HH_DISPLAY_TOPIC 0x0000
#define HH_HELP_FINDER 0x0000
#define HH_DISPLAY_TOC 0x0001
#define HH_DISPLAY_INDEX 0x0002
#define HH_DISPLAY_SEARCH 0x0003
#define HH_SET_WIN_TYPE 0x0004
#define HH_GET_WIN_TYPE 0x0005
#define HH_GET_WIN_HANDLE 0x0006
#define HH_ENUM_INFO_TYPE 0x0007
#define HH_SET_INFO_TYPE 0x0008
#define HH_SYNC 0x0009
#define HH_RESERVED1 0x000A
#define HH_RESERVED2 0x000B
#define HH_RESERVED3 0x000C
#define HH_KEYWORD_LOOKUP 0x000D
#define HH_DISPLAY_TEXT_POPUP 0x000E
#define HH_HELP_CONTEXT 0x000F
#define HH_TP_HELP_CONTEXTMENU 0x0010
#define HH_TP_HELP_WM_HELP 0x0011
#define HH_CLOSE_ALL 0x0012
#define HH_ALINK_LOOKUP 0x0013
#define HH_GET_LAST_ERROR 0x0014
#define HH_ENUM_CATEGORY 0x0015
#define HH_ENUM_CATEGORY_IT 0x0016
#define HH_RESET_IT_FILTER 0x0017
#define HH_SET_INCLUSIVE_FILTER 0x0018
#define HH_SET_EXCLUSIVE_FILTER 0x0019
#define HH_INITIALIZE 0x001C
#define HH_UNINITIALIZE 0x001D
#define HH_PRETRANSLATEMESSAGE 0x00fd
#define HH_SET_GLOBAL_PROPERTY 0x00fc
#define LZERROR_BADINHANDLE (-1)
#define LZERROR_BADOUTHANDLE (-2)
#define LZERROR_READ (-3)
#define LZERROR_WRITE (-4)
#define LZERROR_GLOBALLOC (-5)
#define LZERROR_GLOBLOCK (-6)
#define LZERROR_BADVALUE (-7)
#define LZERROR_UNKNOWNALG (-8)
#define MCIWNDOPENF_NEW 0x0001
#define MCIWNDF_NOAUTOSIZEWINDOW 0x0001
#define MCIWNDF_NOPLAYBAR 0x0002
#define MCIWNDF_NOAUTOSIZEMOVIE 0x0004
#define MCIWNDF_NOMENU 0x0008
#define MCIWNDF_SHOWNAME 0x0010
#define MCIWNDF_SHOWPOS 0x0020
#define MCIWNDF_SHOWMODE 0x0040
#define MCIWNDF_SHOWALL 0x0070
#define MCIWNDF_NOTIFYMODE 0x0100
#define MCIWNDF_NOTIFYPOS 0x0200
#define MCIWNDF_NOTIFYSIZE 0x0400
#define MCIWNDF_NOTIFYERROR 0x1000
#define MCIWNDF_NOTIFYALL 0x1F00
#define MCIWNDF_NOTIFYANSI 0x0080
#define MCIWNDF_NOTIFYMEDIA 0x0880
#define MCIWNDF_RECORD 0x2000
#define MCIWNDF_NOERRORDLG 0x4000
#define MCIWNDF_NOOPEN 0x8000
#define MCIWNDM_GETDEVICEID (WM_USER + 100)
#define MCIWNDM_GETSTART (WM_USER + 103)
#define MCIWNDM_GETLENGTH (WM_USER + 104)
#define MCIWNDM_GETEND (WM_USER + 105)
#define MCIWNDM_EJECT (WM_USER + 107)
#define MCIWNDM_SETZOOM (WM_USER + 108)
#define MCIWNDM_GETZOOM (WM_USER + 109)
#define MCIWNDM_SETVOLUME (WM_USER + 110)
#define MCIWNDM_GETVOLUME (WM_USER + 111)
#define MCIWNDM_SETSPEED (WM_USER + 112)
#define MCIWNDM_GETSPEED (WM_USER + 113)
#define MCIWNDM_SETREPEAT (WM_USER + 114)
#define MCIWNDM_GETREPEAT (WM_USER + 115)
#define MCIWNDM_REALIZE (WM_USER + 118)
#define MCIWNDM_VALIDATEMEDIA (WM_USER + 121)
#define MCIWNDM_PLAYFROM (WM_USER + 122)
#define MCIWNDM_PLAYTO (WM_USER + 123)
#define MCIWNDM_GETPALETTE (WM_USER + 126)
#define MCIWNDM_SETPALETTE (WM_USER + 127)
#define MCIWNDM_SETTIMERS (WM_USER + 129)
#define MCIWNDM_SETACTIVETIMER (WM_USER + 130)
#define MCIWNDM_SETINACTIVETIMER (WM_USER + 131)
#define MCIWNDM_GETACTIVETIMER (WM_USER + 132)
#define MCIWNDM_GETINACTIVETIMER (WM_USER + 133)
#define MCIWNDM_CHANGESTYLES (WM_USER + 135)
#define MCIWNDM_GETSTYLES (WM_USER + 136)
#define MCIWNDM_GETALIAS (WM_USER + 137)
#define MCIWNDM_PLAYREVERSE (WM_USER + 139)
#define MCIWNDM_GET_SOURCE (WM_USER + 140)
#define MCIWNDM_PUT_SOURCE (WM_USER + 141)
#define MCIWNDM_GET_DEST (WM_USER + 142)
#define MCIWNDM_PUT_DEST (WM_USER + 143)
#define MCIWNDM_CAN_PLAY (WM_USER + 144)
#define MCIWNDM_CAN_WINDOW (WM_USER + 145)
#define MCIWNDM_CAN_RECORD (WM_USER + 146)
#define MCIWNDM_CAN_SAVE (WM_USER + 147)
#define MCIWNDM_CAN_EJECT (WM_USER + 148)
#define MCIWNDM_CAN_CONFIG (WM_USER + 149)
#define MCIWNDM_PALETTEKICK (WM_USER + 150)
#define MCIWNDM_OPENINTERFACE (WM_USER + 151)
#define MCIWNDM_SETOWNER (WM_USER + 152)
#define MCIWNDM_SENDSTRING (WM_USER + 101)
#define MCIWNDM_GETPOSITION (WM_USER + 102)
#define MCIWNDM_GETMODE (WM_USER + 106)
#define MCIWNDM_SETTIMEFORMAT (WM_USER + 119)
#define MCIWNDM_GETTIMEFORMAT (WM_USER + 120)
#define MCIWNDM_GETFILENAME (WM_USER + 124)
#define MCIWNDM_GETDEVICE (WM_USER + 125)
#define MCIWNDM_GETERROR (WM_USER + 128)
#define MCIWNDM_NEW (WM_USER + 134)
#define MCIWNDM_RETURNSTRING (WM_USER + 138)
#define MCIWNDM_OPEN (WM_USER + 153)
#define MCIWNDM_NOTIFYMODE (WM_USER + 200)
#define MCIWNDM_NOTIFYPOS (WM_USER + 201)
#define MCIWNDM_NOTIFYSIZE (WM_USER + 202)
#define MCIWNDM_NOTIFYMEDIA (WM_USER + 203)
#define MCIWNDM_NOTIFYERROR (WM_USER + 205)
#define MCIWND_START -1
#define MCIWND_END -2
#define MAXPNAMELEN 32
#define MAXERRORLENGTH 256
#define MAX_JOYSTICKOEMVXDNAME 260
#define MM_MICROSOFT 1
#define MM_MIDI_MAPPER 1
#define MM_WAVE_MAPPER 2
#define MM_SNDBLST_MIDIOUT 3
#define MM_SNDBLST_MIDIIN 4
#define MM_SNDBLST_SYNTH 5
#define MM_SNDBLST_WAVEOUT 6
#define MM_SNDBLST_WAVEIN 7
#define MM_ADLIB 9
#define MM_MPU401_MIDIOUT 10
#define MM_MPU401_MIDIIN 11
#define MM_PC_JOYSTICK 12
#define TIME_MS 0x0001
#define TIME_SAMPLES 0x0002
#define TIME_BYTES 0x0004
#define TIME_SMPTE 0x0008
#define TIME_MIDI 0x0010
#define TIME_TICKS 0x0020
#define MM_JOY1MOVE 0x3A0
#define MM_JOY2MOVE 0x3A1
#define MM_JOY1ZMOVE 0x3A2
#define MM_JOY2ZMOVE 0x3A3
#define MM_JOY1BUTTONDOWN 0x3B5
#define MM_JOY2BUTTONDOWN 0x3B6
#define MM_JOY1BUTTONUP 0x3B7
#define MM_JOY2BUTTONUP 0x3B8
#define MM_MCINOTIFY 0x3B9
#define MM_WOM_OPEN 0x3BB
#define MM_WOM_CLOSE 0x3BC
#define MM_WOM_DONE 0x3BD
#define MM_WIM_OPEN 0x3BE
#define MM_WIM_CLOSE 0x3BF
#define MM_WIM_DATA 0x3C0
#define MM_MIM_OPEN 0x3C1
#define MM_MIM_CLOSE 0x3C2
#define MM_MIM_DATA 0x3C3
#define MM_MIM_LONGDATA 0x3C4
#define MM_MIM_ERROR 0x3C5
#define MM_MIM_LONGERROR 0x3C6
#define MM_MOM_OPEN 0x3C7
#define MM_MOM_CLOSE 0x3C8
#define MM_MOM_DONE 0x3C9
#define MM_DRVM_OPEN 0x3D0
#define MM_DRVM_CLOSE 0x3D1
#define MM_DRVM_DATA 0x3D2
#define MM_DRVM_ERROR 0x3D3
#define MM_STREAM_OPEN 0x3D4
#define MM_STREAM_CLOSE 0x3D5
#define MM_STREAM_DONE 0x3D6
#define MM_STREAM_ERROR 0x3D7
#define MM_MOM_POSITIONCB 0x3CA
#define MM_MCISIGNAL 0x3CB
#define MM_MIM_MOREDATA 0x3CC
#define MM_MIXM_LINE_CHANGE 0x3D0
#define MM_MIXM_CONTROL_CHANGE 0x3D1
#define MMSYSERR_BASE 0
#define WAVERR_BASE 32
#define MIDIERR_BASE 64
#define TIMERR_BASE 96
#define JOYERR_BASE 160
#define MCIERR_BASE 256
#define MIXERR_BASE 1024
#define MCI_STRING_OFFSET 512
#define MCI_VD_OFFSET 1024
#define MCI_CD_OFFSET 1088
#define MCI_WAVE_OFFSET 1152
#define MCI_SEQ_OFFSET 1216
#define MMSYSERR_NOERROR 0
#define MMSYSERR_ERROR (MMSYSERR_BASE + 1)
#define MMSYSERR_BADDEVICEID (MMSYSERR_BASE + 2)
#define MMSYSERR_NOTENABLED (MMSYSERR_BASE + 3)
#define MMSYSERR_ALLOCATED (MMSYSERR_BASE + 4)
#define MMSYSERR_INVALHANDLE (MMSYSERR_BASE + 5)
#define MMSYSERR_NODRIVER (MMSYSERR_BASE + 6)
#define MMSYSERR_NOMEM (MMSYSERR_BASE + 7)
#define MMSYSERR_NOTSUPPORTED (MMSYSERR_BASE + 8)
#define MMSYSERR_BADERRNUM (MMSYSERR_BASE + 9)
#define MMSYSERR_INVALFLAG (MMSYSERR_BASE + 10)
#define MMSYSERR_INVALPARAM (MMSYSERR_BASE + 11)
#define MMSYSERR_HANDLEBUSY (MMSYSERR_BASE + 12)
#define MMSYSERR_INVALIDALIAS (MMSYSERR_BASE + 13)
#define MMSYSERR_BADDB (MMSYSERR_BASE + 14)
#define MMSYSERR_KEYNOTFOUND (MMSYSERR_BASE + 15)
#define MMSYSERR_READERROR (MMSYSERR_BASE + 16)
#define MMSYSERR_WRITEERROR (MMSYSERR_BASE + 17)
#define MMSYSERR_DELETEERROR (MMSYSERR_BASE + 18)
#define MMSYSERR_VALNOTFOUND (MMSYSERR_BASE + 19)
#define MMSYSERR_NODRIVERCB (MMSYSERR_BASE + 20)
#define MMSYSERR_LASTERROR (MMSYSERR_BASE + 20)
#define DRV_LOAD 0x0001
#define DRV_ENABLE 0x0002
#define DRV_OPEN 0x0003
#define DRV_CLOSE 0x0004
#define DRV_DISABLE 0x0005
#define DRV_FREE 0x0006
#define DRV_CONFIGURE 0x0007
#define DRV_QUERYCONFIGURE 0x0008
#define DRV_INSTALL 0x0009
#define DRV_REMOVE 0x000A
#define DRV_EXITSESSION 0x000B
#define DRV_POWER 0x000F
#define DRV_RESERVED 0x0800
#define DRV_USER 0x4000
#define DRVCNF_CANCEL 0x0000
#define DRVCNF_OK 0x0001
#define DRVCNF_RESTART 0x0002
#define DRV_CANCEL DRVCNF_CANCEL
#define DRV_OK DRVCNF_OK
#define DRV_RESTART DRVCNF_RESTART
#define DRV_MCI_FIRST DRV_RESERVED
#define DRV_MCI_LAST (DRV_RESERVED + 0xFFF)
#define CALLBACK_TYPEMASK 0x00070000l
#define CALLBACK_NULL 0x00000000l
#define CALLBACK_WINDOW 0x00010000l
#define CALLBACK_TASK 0x00020000l
#define CALLBACK_FUNCTION 0x00030000l
#define CALLBACK_THREAD (CALLBACK_TASK)
#define CALLBACK_EVENT 0x00050000l
#define SND_SYNC 0x0000
#define SND_ASYNC 0x0001
#define SND_NODEFAULT 0x0002
#define SND_MEMORY 0x0004
#define SND_LOOP 0x0008
#define SND_NOSTOP 0x0010
#define SND_NOWAIT 0x00002000L
#define SND_ALIAS 0x00010000L
#define SND_ALIAS_ID 0x00110000L
#define SND_FILENAME 0x00020000L
#define SND_RESOURCE 0x00040004L
#define SND_PURGE 0x0040
#define SND_APPLICATION 0x0080
#define SND_ALIAS_START 0
#define WAVERR_BADFORMAT (WAVERR_BASE + 0)
#define WAVERR_STILLPLAYING (WAVERR_BASE + 1)
#define WAVERR_UNPREPARED (WAVERR_BASE + 2)
#define WAVERR_SYNC (WAVERR_BASE + 3)
#define WAVERR_LASTERROR (WAVERR_BASE + 3)
#define WOM_OPEN MM_WOM_OPEN
#define WOM_CLOSE MM_WOM_CLOSE
#define WOM_DONE MM_WOM_DONE
#define WIM_OPEN MM_WIM_OPEN
#define WIM_CLOSE MM_WIM_CLOSE
#define WIM_DATA MM_WIM_DATA
#define WAVE_MAPPER -1
#define WAVE_FORMAT_QUERY 0x0001
#define WAVE_ALLOWSYNC 0x0002
#define WAVE_MAPPED 0x0004
#define WHDR_DONE 0x00000001
#define WHDR_PREPARED 0x00000002
#define WHDR_BEGINLOOP 0x00000004
#define WHDR_ENDLOOP 0x00000008
#define WHDR_INQUEUE 0x00000010
#define WAVECAPS_PITCH 0x0001
#define WAVECAPS_PLAYBACKRATE 0x0002
#define WAVECAPS_VOLUME 0x0004
#define WAVECAPS_LRVOLUME 0x0008
#define WAVECAPS_SYNC 0x0010
#define WAVECAPS_SAMPLEACCURATE 0x0020
#define WAVECAPS_DIRECTSOUND 0x0040
#define WAVE_INVALIDFORMAT 0x00000000
#define WAVE_FORMAT_1M08 0x00000001
#define WAVE_FORMAT_1S08 0x00000002
#define WAVE_FORMAT_1M16 0x00000004
#define WAVE_FORMAT_1S16 0x00000008
#define WAVE_FORMAT_2M08 0x00000010
#define WAVE_FORMAT_2S08 0x00000020
#define WAVE_FORMAT_2M16 0x00000040
#define WAVE_FORMAT_2S16 0x00000080
#define WAVE_FORMAT_4M08 0x00000100
#define WAVE_FORMAT_4S08 0x00000200
#define WAVE_FORMAT_4M16 0x00000400
#define WAVE_FORMAT_4S16 0x00000800
#define WAVE_FORMAT_PCM 1
#define MIDIERR_UNPREPARED (MIDIERR_BASE + 0)
#define MIDIERR_STILLPLAYING (MIDIERR_BASE + 1)
#define MIDIERR_NOMAP (MIDIERR_BASE + 2)
#define MIDIERR_NOTREADY (MIDIERR_BASE + 3)
#define MIDIERR_NODEVICE (MIDIERR_BASE + 4)
#define MIDIERR_INVALIDSETUP (MIDIERR_BASE + 5)
#define MIDIERR_BADOPENMODE (MIDIERR_BASE + 6)
#define MIDIERR_DONT_CONTINUE (MIDIERR_BASE + 7)
#define MIDIERR_LASTERROR (MIDIERR_BASE + 7)
#define MIDIPATCHSIZE 128
#define MIM_OPEN MM_MIM_OPEN
#define MIM_CLOSE MM_MIM_CLOSE
#define MIM_DATA MM_MIM_DATA
#define MIM_LONGDATA MM_MIM_LONGDATA
#define MIM_ERROR MM_MIM_ERROR
#define MIM_LONGERROR MM_MIM_LONGERROR
#define MOM_OPEN MM_MOM_OPEN
#define MOM_CLOSE MM_MOM_CLOSE
#define MOM_DONE MM_MOM_DONE
#define MIM_MOREDATA MM_MIM_MOREDATA
#define MOM_POSITIONCB MM_MOM_POSITIONCB
#define MIDIMAPPER -1
#define MIDI_MAPPER -1
#define MIDI_IO_STATUS 0x00000020L
#define MIDI_CACHE_ALL 1
#define MIDI_CACHE_BESTFIT 2
#define MIDI_CACHE_QUERY 3
#define MIDI_UNCACHE 4
#define MOD_MIDIPORT 1
#define MOD_SYNTH 2
#define MOD_SQSYNTH 3
#define MOD_FMSYNTH 4
#define MOD_MAPPER 5
#define MIDICAPS_VOLUME 0x0001
#define MIDICAPS_LRVOLUME 0x0002
#define MIDICAPS_CACHE 0x0004
#define MIDICAPS_STREAM 0x0008
#define MHDR_DONE 0x00000001
#define MHDR_PREPARED 0x00000002
#define MHDR_INQUEUE 0x00000004
#define MHDR_ISSTRM 0x00000008
#define MEVT_F_SHORT 0x00000000L
#define MEVT_F_LONG 0x80000000L
#define MEVT_F_CALLBACK 0x40000000L
#define MEVT_SHORTMSG BYTE(_CAST, 0x00)
#define MEVT_TEMPO BYTE(_CAST, 0x01)
#define MEVT_NOP BYTE(_CAST, 0x02)
#define MEVT_LONGMSG BYTE(_CAST, 0x80)
#define MEVT_COMMENT BYTE(_CAST, 0x82)
#define MEVT_VERSION BYTE(_CAST, 0x84)
#define MIDISTRM_ERROR (-2)
#define MIDIPROP_SET 0x80000000L
#define MIDIPROP_GET 0x40000000L
#define MIDIPROP_TIMEDIV 0x00000001L
#define MIDIPROP_TEMPO 0x00000002L
#define AUX_MAPPER -1
#define AUXCAPS_CDAUDIO 1
#define AUXCAPS_AUXIN 2
#define AUXCAPS_VOLUME 0x0001
#define AUXCAPS_LRVOLUME 0x0002
#define MIXER_SHORT_NAME_CHARS 16
#define MIXER_LONG_NAME_CHARS 64
#define MIXERR_INVALLINE (MIXERR_BASE + 0)
#define MIXERR_INVALCONTROL (MIXERR_BASE + 1)
#define MIXERR_INVALVALUE (MIXERR_BASE + 2)
#define MIXERR_LASTERROR (MIXERR_BASE + 2)
#define MIXER_OBJECTF_HANDLE 0x80000000L
#define MIXER_OBJECTF_MIXER 0x00000000L
#define MIXER_OBJECTF_HMIXER 0x80000000L
#define MIXER_OBJECTF_WAVEOUT 0x10000000L
#define MIXER_OBJECTF_HWAVEOUT 0x90000000L
#define MIXER_OBJECTF_WAVEIN 0x20000000L
#define MIXER_OBJECTF_HWAVEIN 0xA0000000L
#define MIXER_OBJECTF_MIDIOUT 0x30000000L
#define MIXER_OBJECTF_HMIDIOUT 0xB0000000L
#define MIXER_OBJECTF_MIDIIN 0x40000000L
#define MIXER_OBJECTF_HMIDIIN 0xC0000000L
#define MIXER_OBJECTF_AUX 0x50000000L
#define MIXERLINE_LINEF_ACTIVE 0x00000001L
#define MIXERLINE_LINEF_DISCONNECTED 0x00008000L
#define MIXERLINE_LINEF_SOURCE 0x80000000L
#define MIXERLINE_COMPONENTTYPE_DST_FIRST 0x00000000L
#define MIXERLINE_COMPONENTTYPE_DST_UNDEFINED (MIXERLINE_COMPONENTTYPE_DST_FIRST + 0)
#define MIXERLINE_COMPONENTTYPE_DST_DIGITAL (MIXERLINE_COMPONENTTYPE_DST_FIRST + 1)
#define MIXERLINE_COMPONENTTYPE_DST_LINE (MIXERLINE_COMPONENTTYPE_DST_FIRST + 2)
#define MIXERLINE_COMPONENTTYPE_DST_MONITOR (MIXERLINE_COMPONENTTYPE_DST_FIRST + 3)
#define MIXERLINE_COMPONENTTYPE_DST_SPEAKERS (MIXERLINE_COMPONENTTYPE_DST_FIRST + 4)
#define MIXERLINE_COMPONENTTYPE_DST_HEADPHONES (MIXERLINE_COMPONENTTYPE_DST_FIRST + 5)
#define MIXERLINE_COMPONENTTYPE_DST_TELEPHONE (MIXERLINE_COMPONENTTYPE_DST_FIRST + 6)
#define MIXERLINE_COMPONENTTYPE_DST_WAVEIN (MIXERLINE_COMPONENTTYPE_DST_FIRST + 7)
#define MIXERLINE_COMPONENTTYPE_DST_VOICEIN (MIXERLINE_COMPONENTTYPE_DST_FIRST + 8)
#define MIXERLINE_COMPONENTTYPE_DST_LAST (MIXERLINE_COMPONENTTYPE_DST_FIRST + 8)
#define MIXERLINE_COMPONENTTYPE_SRC_FIRST 0x00001000L
#define MIXERLINE_COMPONENTTYPE_SRC_UNDEFINED (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 0)
#define MIXERLINE_COMPONENTTYPE_SRC_DIGITAL (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 1)
#define MIXERLINE_COMPONENTTYPE_SRC_LINE (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 2)
#define MIXERLINE_COMPONENTTYPE_SRC_MICROPHONE (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 3)
#define MIXERLINE_COMPONENTTYPE_SRC_SYNTHESIZER (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 4)
#define MIXERLINE_COMPONENTTYPE_SRC_COMPACTDISC (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 5)
#define MIXERLINE_COMPONENTTYPE_SRC_TELEPHONE (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 6)
#define MIXERLINE_COMPONENTTYPE_SRC_PCSPEAKER (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 7)
#define MIXERLINE_COMPONENTTYPE_SRC_WAVEOUT (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 8)
#define MIXERLINE_COMPONENTTYPE_SRC_AUXILIARY (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 9)
#define MIXERLINE_COMPONENTTYPE_SRC_ANALOG (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 10)
#define MIXERLINE_COMPONENTTYPE_SRC_LAST (MIXERLINE_COMPONENTTYPE_SRC_FIRST + 10)
#define MIXERLINE_TARGETTYPE_UNDEFINED 0
#define MIXERLINE_TARGETTYPE_WAVEOUT 1
#define MIXERLINE_TARGETTYPE_WAVEIN 2
#define MIXERLINE_TARGETTYPE_MIDIOUT 3
#define MIXERLINE_TARGETTYPE_MIDIIN 4
#define MIXERLINE_TARGETTYPE_AUX 5
#define MIXER_GETLINEINFOF_DESTINATION 0x00000000L
#define MIXER_GETLINEINFOF_SOURCE 0x00000001L
#define MIXER_GETLINEINFOF_LINEID 0x00000002L
#define MIXER_GETLINEINFOF_COMPONENTTYPE 0x00000003L
#define MIXER_GETLINEINFOF_TARGETTYPE 0x00000004L
#define MIXER_GETLINEINFOF_QUERYMASK 0x0000000FL
#define MIXERCONTROL_CONTROLF_UNIFORM 0x00000001L
#define MIXERCONTROL_CONTROLF_MULTIPLE 0x00000002L
#define MIXERCONTROL_CONTROLF_DISABLED 0x80000000L
#define MIXERCONTROL_CT_CLASS_MASK 0xF0000000L
#define MIXERCONTROL_CT_CLASS_CUSTOM 0x00000000L
#define MIXERCONTROL_CT_CLASS_METER 0x10000000L
#define MIXERCONTROL_CT_CLASS_SWITCH 0x20000000L
#define MIXERCONTROL_CT_CLASS_NUMBER 0x30000000L
#define MIXERCONTROL_CT_CLASS_SLIDER 0x40000000L
#define MIXERCONTROL_CT_CLASS_FADER 0x50000000L
#define MIXERCONTROL_CT_CLASS_TIME 0x60000000L
#define MIXERCONTROL_CT_CLASS_LIST 0x70000000L
#define MIXERCONTROL_CT_SUBCLASS_MASK 0x0F000000L
#define MIXERCONTROL_CT_SC_SWITCH_BOOLEAN 0x00000000L
#define MIXERCONTROL_CT_SC_SWITCH_BUTTON 0x01000000L
#define MIXERCONTROL_CT_SC_METER_POLLED 0x00000000L
#define MIXERCONTROL_CT_SC_TIME_MICROSECS 0x00000000L
#define MIXERCONTROL_CT_SC_TIME_MILLISECS 0x01000000L
#define MIXERCONTROL_CT_SC_LIST_SINGLE 0x00000000L
#define MIXERCONTROL_CT_SC_LIST_MULTIPLE 0x01000000L
#define MIXERCONTROL_CT_UNITS_MASK 0x00FF0000L
#define MIXERCONTROL_CT_UNITS_CUSTOM 0x00000000L
#define MIXERCONTROL_CT_UNITS_BOOLEAN 0x00010000L
#define MIXERCONTROL_CT_UNITS_SIGNED 0x00020000L
#define MIXERCONTROL_CT_UNITS_UNSIGNED 0x00030000L
#define MIXERCONTROL_CT_UNITS_DECIBELS 0x00040000L
#define MIXERCONTROL_CT_UNITS_PERCENT 0x00050000L
#define MIXERCONTROL_CONTROLTYPE_CUSTOM 0x00000000L
#define MIXERCONTROL_CONTROLTYPE_BOOLEANMETER 0x10010000L
#define MIXERCONTROL_CONTROLTYPE_SIGNEDMETER 0x10020000L
#define MIXERCONTROL_CONTROLTYPE_PEAKMETER (MIXERCONTROL_CONTROLTYPE_SIGNEDMETER + 1)
#define MIXERCONTROL_CONTROLTYPE_UNSIGNEDMETER 0x10030000L
#define MIXERCONTROL_CONTROLTYPE_BOOLEAN 0x20010000L
#define MIXERCONTROL_CONTROLTYPE_ONOFF (MIXERCONTROL_CONTROLTYPE_BOOLEAN + 1)
#define MIXERCONTROL_CONTROLTYPE_MUTE (MIXERCONTROL_CONTROLTYPE_BOOLEAN + 2)
#define MIXERCONTROL_CONTROLTYPE_MONO (MIXERCONTROL_CONTROLTYPE_BOOLEAN + 3)
#define MIXERCONTROL_CONTROLTYPE_LOUDNESS (MIXERCONTROL_CONTROLTYPE_BOOLEAN + 4)
#define MIXERCONTROL_CONTROLTYPE_STEREOENH (MIXERCONTROL_CONTROLTYPE_BOOLEAN + 5)
#define MIXERCONTROL_CONTROLTYPE_BUTTON 0x21010000L
#define MIXERCONTROL_CONTROLTYPE_DECIBELS 0x30040000L
#define MIXERCONTROL_CONTROLTYPE_SIGNED 0x30020000L
#define MIXERCONTROL_CONTROLTYPE_UNSIGNED 0x30030000L
#define MIXERCONTROL_CONTROLTYPE_PERCENT 0x30050000L
#define MIXERCONTROL_CONTROLTYPE_SLIDER 0x40020000L
#define MIXERCONTROL_CONTROLTYPE_PAN (MIXERCONTROL_CONTROLTYPE_SLIDER + 1)
#define MIXERCONTROL_CONTROLTYPE_QSOUNDPAN (MIXERCONTROL_CONTROLTYPE_SLIDER + 2)
#define MIXERCONTROL_CONTROLTYPE_FADER 0x50030000L
#define MIXERCONTROL_CONTROLTYPE_VOLUME (MIXERCONTROL_CONTROLTYPE_FADER + 1)
#define MIXERCONTROL_CONTROLTYPE_BASS (MIXERCONTROL_CONTROLTYPE_FADER + 2)
#define MIXERCONTROL_CONTROLTYPE_TREBLE (MIXERCONTROL_CONTROLTYPE_FADER + 3)
#define MIXERCONTROL_CONTROLTYPE_EQUALIZER (MIXERCONTROL_CONTROLTYPE_FADER + 4)
#define MIXERCONTROL_CONTROLTYPE_SINGLESELECT 0x70010000L
#define MIXERCONTROL_CONTROLTYPE_MUX (MIXERCONTROL_CONTROLTYPE_SINGLESELECT + 1)
#define MIXERCONTROL_CONTROLTYPE_MULTIPLESELECT 0x71010000L
#define MIXERCONTROL_CONTROLTYPE_MIXER (MIXERCONTROL_CONTROLTYPE_MULTIPLESELECT + 1)
#define MIXERCONTROL_CONTROLTYPE_MICROTIME 0x60030000L
#define MIXERCONTROL_CONTROLTYPE_MILLITIME 0x61030000L
#define MIXER_GETLINECONTROLSF_ALL 0x00000000L
#define MIXER_GETLINECONTROLSF_ONEBYID 0x00000001L
#define MIXER_GETLINECONTROLSF_ONEBYTYPE 0x00000002L
#define MIXER_GETLINECONTROLSF_QUERYMASK 0x0000000FL
#define MIXER_GETCONTROLDETAILSF_VALUE 0x00000000L
#define MIXER_GETCONTROLDETAILSF_LISTTEXT 0x00000001L
#define MIXER_GETCONTROLDETAILSF_QUERYMASK 0x0000000FL
#define MIXER_SETCONTROLDETAILSF_VALUE 0x00000000L
#define MIXER_SETCONTROLDETAILSF_CUSTOM 0x00000001L
#define MIXER_SETCONTROLDETAILSF_QUERYMASK 0x0000000FL
#define TIMERR_NOERROR (0)
#define TIMERR_NOCANDO (TIMERR_BASE+1)
#define TIMERR_STRUCT (TIMERR_BASE+33)
#define TIME_ONESHOT 0x0000
#define TIME_PERIODIC 0x0001
#define TIME_CALLBACK_FUNCTION 0x0000
#define TIME_CALLBACK_EVENT_SET 0x0010
#define TIME_CALLBACK_EVENT_PULSE 0x0020
#define JOYERR_NOERROR (0)
#define JOYERR_PARMS (JOYERR_BASE+5)
#define JOYERR_NOCANDO (JOYERR_BASE+6)
#define JOYERR_UNPLUGGED (JOYERR_BASE+7)
#define JOY_BUTTON1 0x0001
#define JOY_BUTTON2 0x0002
#define JOY_BUTTON3 0x0004
#define JOY_BUTTON4 0x0008
#define JOY_BUTTON1CHG 0x0100
#define JOY_BUTTON2CHG 0x0200
#define JOY_BUTTON3CHG 0x0400
#define JOY_BUTTON4CHG 0x0800
#define JOY_BUTTON5 0x00000010l
#define JOY_BUTTON6 0x00000020l
#define JOY_BUTTON7 0x00000040l
#define JOY_BUTTON8 0x00000080l
#define JOY_BUTTON9 0x00000100l
#define JOY_BUTTON10 0x00000200l
#define JOY_BUTTON11 0x00000400l
#define JOY_BUTTON12 0x00000800l
#define JOY_BUTTON13 0x00001000l
#define JOY_BUTTON14 0x00002000l
#define JOY_BUTTON15 0x00004000l
#define JOY_BUTTON16 0x00008000l
#define JOY_BUTTON17 0x00010000l
#define JOY_BUTTON18 0x00020000l
#define JOY_BUTTON19 0x00040000l
#define JOY_BUTTON20 0x00080000l
#define JOY_BUTTON21 0x00100000l
#define JOY_BUTTON22 0x00200000l
#define JOY_BUTTON23 0x00400000l
#define JOY_BUTTON24 0x00800000l
#define JOY_BUTTON25 0x01000000l
#define JOY_BUTTON26 0x02000000l
#define JOY_BUTTON27 0x04000000l
#define JOY_BUTTON28 0x08000000l
#define JOY_BUTTON29 0x10000000l
#define JOY_BUTTON30 0x20000000l
#define JOY_BUTTON31 0x40000000l
#define JOY_BUTTON32 0x80000000l
#define JOY_POVCENTERED -1
#define JOY_POVFORWARD 0
#define JOY_POVRIGHT 9000
#define JOY_POVBACKWARD 18000
#define JOY_POVLEFT 27000
#define JOY_RETURNX 0x00000001l
#define JOY_RETURNY 0x00000002l
#define JOY_RETURNZ 0x00000004l
#define JOY_RETURNR 0x00000008l
#define JOY_RETURNU 0x00000010l
#define JOY_RETURNV 0x00000020l
#define JOY_RETURNPOV 0x00000040l
#define JOY_RETURNBUTTONS 0x00000080l
#define JOY_RETURNRAWDATA 0x00000100l
#define JOY_RETURNPOVCTS 0x00000200l
#define JOY_RETURNCENTERED 0x00000400l
#define JOY_USEDEADZONE 0x00000800l
#define JOY_RETURNALL 0x000000FFl
#define JOY_CAL_READALWAYS 0x00010000l
#define JOY_CAL_READXYONLY 0x00020000l
#define JOY_CAL_READ3 0x00040000l
#define JOY_CAL_READ4 0x00080000l
#define JOY_CAL_READXONLY 0x00100000l
#define JOY_CAL_READYONLY 0x00200000l
#define JOY_CAL_READ5 0x00400000l
#define JOY_CAL_READ6 0x00800000l
#define JOY_CAL_READZONLY 0x01000000l
#define JOY_CAL_READRONLY 0x02000000l
#define JOY_CAL_READUONLY 0x04000000l
#define JOY_CAL_READVONLY 0x08000000l
#define JOYSTICKID1 0
#define JOYSTICKID2 1
#define JOYCAPS_HASZ 0x0001
#define JOYCAPS_HASR 0x0002
#define JOYCAPS_HASU 0x0004
#define JOYCAPS_HASV 0x0008
#define JOYCAPS_HASPOV 0x0010
#define JOYCAPS_POV4DIR 0x0020
#define JOYCAPS_POVCTS 0x0040
#define MMIOERR_BASE 256
#define MMIOERR_FILENOTFOUND (MMIOERR_BASE + 1)
#define MMIOERR_OUTOFMEMORY (MMIOERR_BASE + 2)
#define MMIOERR_CANNOTOPEN (MMIOERR_BASE + 3)
#define MMIOERR_CANNOTCLOSE (MMIOERR_BASE + 4)
#define MMIOERR_CANNOTREAD (MMIOERR_BASE + 5)
#define MMIOERR_CANNOTWRITE (MMIOERR_BASE + 6)
#define MMIOERR_CANNOTSEEK (MMIOERR_BASE + 7)
#define MMIOERR_CANNOTEXPAND (MMIOERR_BASE + 8)
#define MMIOERR_CHUNKNOTFOUND (MMIOERR_BASE + 9)
#define MMIOERR_UNBUFFERED (MMIOERR_BASE + 10)
#define MMIOERR_PATHNOTFOUND (MMIOERR_BASE + 11)
#define MMIOERR_ACCESSDENIED (MMIOERR_BASE + 12)
#define MMIOERR_SHARINGVIOLATION (MMIOERR_BASE + 13)
#define MMIOERR_NETWORKERROR (MMIOERR_BASE + 14)
#define MMIOERR_TOOMANYOPENFILES (MMIOERR_BASE + 15)
#define MMIOERR_INVALIDFILE (MMIOERR_BASE + 16)
#define CFSEPCHAR "+"
#define MMIO_RWMODE 0x00000003
#define MMIO_SHAREMODE 0x00000070
#define MMIO_CREATE 0x00001000
#define MMIO_PARSE 0x00000100
#define MMIO_DELETE 0x00000200
#define MMIO_EXIST 0x00004000
#define MMIO_ALLOCBUF 0x00010000
#define MMIO_GETTEMP 0x00020000
#define MMIO_DIRTY 0x10000000
#define MMIO_READ 0x00000000
#define MMIO_WRITE 0x00000001
#define MMIO_READWRITE 0x00000002
#define MMIO_COMPAT 0x00000000
#define MMIO_EXCLUSIVE 0x00000010
#define MMIO_DENYWRITE 0x00000020
#define MMIO_DENYREAD 0x00000030
#define MMIO_DENYNONE 0x00000040
#define MMIO_FHOPEN 0x0010
#define MMIO_EMPTYBUF 0x0010
#define MMIO_TOUPPER 0x0010
#define MMIO_INSTALLPROC 0x00010000
#define MMIO_GLOBALPROC 0x10000000
#define MMIO_REMOVEPROC 0x00020000
#define MMIO_UNICODEPROC 0x01000000
#define MMIO_FINDPROC 0x00040000
#define MMIO_FINDCHUNK 0x0010
#define MMIO_FINDRIFF 0x0020
#define MMIO_FINDLIST 0x0040
#define MMIO_CREATERIFF 0x0020
#define MMIO_CREATELIST 0x0040
#define MMIOM_READ MMIO_READ
#define MMIOM_WRITE MMIO_WRITE
#define MMIOM_SEEK 2
#define MMIOM_OPEN 3
#define MMIOM_CLOSE 4
#define MMIOM_WRITEFLUSH 5
#define MMIOM_RENAME 6
#define MMIOM_USER 0x8000
#define FOURCC_RIFF dword(_cast, 0x46464952)
#define FOURCC_LIST dword(_cast, 0x5453494C)
#define FOURCC_DOS dword(_cast, 0x20534F44)
#define FOURCC_MEM dword(_cast, 0x204D454D)
#define SEEK_SET 0
#define SEEK_CUR 1
#define SEEK_END 2
#define MMIO_DEFAULTBUFFER 8192
#define MCIERR_INVALID_DEVICE_ID (MCIERR_BASE + 1)
#define MCIERR_UNRECOGNIZED_KEYWORD (MCIERR_BASE + 3)
#define MCIERR_UNRECOGNIZED_COMMAND (MCIERR_BASE + 5)
#define MCIERR_HARDWARE (MCIERR_BASE + 6)
#define MCIERR_INVALID_DEVICE_NAME (MCIERR_BASE + 7)
#define MCIERR_OUT_OF_MEMORY (MCIERR_BASE + 8)
#define MCIERR_DEVICE_OPEN (MCIERR_BASE + 9)
#define MCIERR_CANNOT_LOAD_DRIVER (MCIERR_BASE + 10)
#define MCIERR_MISSING_COMMAND_STRING (MCIERR_BASE + 11)
#define MCIERR_PARAM_OVERFLOW (MCIERR_BASE + 12)
#define MCIERR_MISSING_STRING_ARGUMENT (MCIERR_BASE + 13)
#define MCIERR_BAD_INTEGER (MCIERR_BASE + 14)
#define MCIERR_PARSER_INTERNAL (MCIERR_BASE + 15)
#define MCIERR_DRIVER_INTERNAL (MCIERR_BASE + 16)
#define MCIERR_MISSING_PARAMETER (MCIERR_BASE + 17)
#define MCIERR_UNSUPPORTED_FUNCTION (MCIERR_BASE + 18)
#define MCIERR_FILE_NOT_FOUND (MCIERR_BASE + 19)
#define MCIERR_DEVICE_NOT_READY (MCIERR_BASE + 20)
#define MCIERR_INTERNAL (MCIERR_BASE + 21)
#define MCIERR_DRIVER (MCIERR_BASE + 22)
#define MCIERR_CANNOT_USE_ALL (MCIERR_BASE + 23)
#define MCIERR_MULTIPLE (MCIERR_BASE + 24)
#define MCIERR_EXTENSION_NOT_FOUND (MCIERR_BASE + 25)
#define MCIERR_OUTOFRANGE (MCIERR_BASE + 26)
#define MCIERR_FLAGS_NOT_COMPATIBLE (MCIERR_BASE + 28)
#define MCIERR_FILE_NOT_SAVED (MCIERR_BASE + 30)
#define MCIERR_DEVICE_TYPE_REQUIRED (MCIERR_BASE + 31)
#define MCIERR_DEVICE_LOCKED (MCIERR_BASE + 32)
#define MCIERR_DUPLICATE_ALIAS (MCIERR_BASE + 33)
#define MCIERR_BAD_CONSTANT (MCIERR_BASE + 34)
#define MCIERR_MUST_USE_SHAREABLE (MCIERR_BASE + 35)
#define MCIERR_MISSING_DEVICE_NAME (MCIERR_BASE + 36)
#define MCIERR_BAD_TIME_FORMAT (MCIERR_BASE + 37)
#define MCIERR_NO_CLOSING_QUOTE (MCIERR_BASE + 38)
#define MCIERR_DUPLICATE_FLAGS (MCIERR_BASE + 39)
#define MCIERR_INVALID_FILE (MCIERR_BASE + 40)
#define MCIERR_NULL_PARAMETER_BLOCK (MCIERR_BASE + 41)
#define MCIERR_UNNAMED_RESOURCE (MCIERR_BASE + 42)
#define MCIERR_NEW_REQUIRES_ALIAS (MCIERR_BASE + 43)
#define MCIERR_NOTIFY_ON_AUTO_OPEN (MCIERR_BASE + 44)
#define MCIERR_NO_ELEMENT_ALLOWED (MCIERR_BASE + 45)
#define MCIERR_NONAPPLICABLE_FUNCTION (MCIERR_BASE + 46)
#define MCIERR_ILLEGAL_FOR_AUTO_OPEN (MCIERR_BASE + 47)
#define MCIERR_FILENAME_REQUIRED (MCIERR_BASE + 48)
#define MCIERR_EXTRA_CHARACTERS (MCIERR_BASE + 49)
#define MCIERR_DEVICE_NOT_INSTALLED (MCIERR_BASE + 50)
#define MCIERR_GET_CD (MCIERR_BASE + 51)
#define MCIERR_SET_CD (MCIERR_BASE + 52)
#define MCIERR_SET_DRIVE (MCIERR_BASE + 53)
#define MCIERR_DEVICE_LENGTH (MCIERR_BASE + 54)
#define MCIERR_DEVICE_ORD_LENGTH (MCIERR_BASE + 55)
#define MCIERR_NO_INTEGER (MCIERR_BASE + 56)
#define MCIERR_WAVE_OUTPUTSINUSE (MCIERR_BASE + 64)
#define MCIERR_WAVE_SETOUTPUTINUSE (MCIERR_BASE + 65)
#define MCIERR_WAVE_INPUTSINUSE (MCIERR_BASE + 66)
#define MCIERR_WAVE_SETINPUTINUSE (MCIERR_BASE + 67)
#define MCIERR_WAVE_OUTPUTUNSPECIFIED (MCIERR_BASE + 68)
#define MCIERR_WAVE_INPUTUNSPECIFIED (MCIERR_BASE + 69)
#define MCIERR_WAVE_OUTPUTSUNSUITABLE (MCIERR_BASE + 70)
#define MCIERR_WAVE_SETOUTPUTUNSUITABLE (MCIERR_BASE + 71)
#define MCIERR_WAVE_INPUTSUNSUITABLE (MCIERR_BASE + 72)
#define MCIERR_WAVE_SETINPUTUNSUITABLE (MCIERR_BASE + 73)
#define MCIERR_SEQ_DIV_INCOMPATIBLE (MCIERR_BASE + 80)
#define MCIERR_SEQ_PORT_INUSE (MCIERR_BASE + 81)
#define MCIERR_SEQ_PORT_NONEXISTENT (MCIERR_BASE + 82)
#define MCIERR_SEQ_PORT_MAPNODEVICE (MCIERR_BASE + 83)
#define MCIERR_SEQ_PORT_MISCERROR (MCIERR_BASE + 84)
#define MCIERR_SEQ_TIMER (MCIERR_BASE + 85)
#define MCIERR_SEQ_PORTUNSPECIFIED (MCIERR_BASE + 86)
#define MCIERR_SEQ_NOMIDIPRESENT (MCIERR_BASE + 87)
#define MCIERR_NO_WINDOW (MCIERR_BASE + 90)
#define MCIERR_CREATEWINDOW (MCIERR_BASE + 91)
#define MCIERR_FILE_READ (MCIERR_BASE + 92)
#define MCIERR_FILE_WRITE (MCIERR_BASE + 93)
#define MCIERR_NO_IDENTITY (MCIERR_BASE + 94)
#define MCIERR_CUSTOM_DRIVER_BASE (MCIERR_BASE + 256)
#define MCI_FIRST DRV_MCI_FIRST
#define MCI_OPEN 0x0803
#define MCI_CLOSE 0x0804
#define MCI_ESCAPE 0x0805
#define MCI_PLAY 0x0806
#define MCI_SEEK 0x0807
#define MCI_STOP 0x0808
#define MCI_PAUSE 0x0809
#define MCI_INFO 0x080A
#define MCI_GETDEVCAPS 0x080B
#define MCI_SPIN 0x080C
#define MCI_SET 0x080D
#define MCI_STEP 0x080E
#define MCI_RECORD 0x080F
#define MCI_SYSINFO 0x0810
#define MCI_BREAK 0x0811
#define MCI_SAVE 0x0813
#define MCI_STATUS 0x0814
#define MCI_CUE 0x0830
#define MCI_REALIZE 0x0840
#define MCI_WINDOW 0x0841
#define MCI_PUT 0x0842
#define MCI_WHERE 0x0843
#define MCI_FREEZE 0x0844
#define MCI_UNFREEZE 0x0845
#define MCI_LOAD 0x0850
#define MCI_CUT 0x0851
#define MCI_COPY 0x0852
#define MCI_PASTE 0x0853
#define MCI_UPDATE 0x0854
#define MCI_RESUME 0x0855
#define MCI_DELETE 0x0856
#define MCI_USER_MESSAGES (DRV_MCI_FIRST + 0x400)
#define MCI_LAST 0x0FFF
#define MCI_ALL_DEVICE_ID -1
#define MCI_DEVTYPE_VCR 513
#define MCI_DEVTYPE_VIDEODISC 514
#define MCI_DEVTYPE_OVERLAY 515
#define MCI_DEVTYPE_CD_AUDIO 516
#define MCI_DEVTYPE_DAT 517
#define MCI_DEVTYPE_SCANNER 518
#define MCI_DEVTYPE_ANIMATION 519
#define MCI_DEVTYPE_DIGITAL_VIDEO 520
#define MCI_DEVTYPE_OTHER 521
#define MCI_DEVTYPE_WAVEFORM_AUDIO 522
#define MCI_DEVTYPE_SEQUENCER 523
#define MCI_DEVTYPE_FIRST MCI_DEVTYPE_VCR
#define MCI_DEVTYPE_LAST MCI_DEVTYPE_SEQUENCER
#define MCI_DEVTYPE_FIRST_USER 0x1000
#define MCI_MODE_NOT_READY (MCI_STRING_OFFSET + 12)
#define MCI_MODE_STOP (MCI_STRING_OFFSET + 13)
#define MCI_MODE_PLAY (MCI_STRING_OFFSET + 14)
#define MCI_MODE_RECORD (MCI_STRING_OFFSET + 15)
#define MCI_MODE_SEEK (MCI_STRING_OFFSET + 16)
#define MCI_MODE_PAUSE (MCI_STRING_OFFSET + 17)
#define MCI_MODE_OPEN (MCI_STRING_OFFSET + 18)
#define MCI_FORMAT_MILLISECONDS 0
#define MCI_FORMAT_HMS 1
#define MCI_FORMAT_MSF 2
#define MCI_FORMAT_FRAMES 3
#define MCI_FORMAT_SMPTE_24 4
#define MCI_FORMAT_SMPTE_25 5
#define MCI_FORMAT_SMPTE_30 6
#define MCI_FORMAT_SMPTE_30DROP 7
#define MCI_FORMAT_BYTES 8
#define MCI_FORMAT_SAMPLES 9
#define MCI_FORMAT_TMSF 10
#define MCI_NOTIFY_SUCCESSFUL 0x0001
#define MCI_NOTIFY_SUPERSEDED 0x0002
#define MCI_NOTIFY_ABORTED 0x0004
#define MCI_NOTIFY_FAILURE 0x0008
#define MCI_NOTIFY 0x00000001L
#define MCI_WAIT 0x00000002L
#define MCI_FROM 0x00000004L
#define MCI_TO 0x00000008L
#define MCI_TRACK 0x00000010L
#define MCI_OPEN_SHAREABLE 0x00000100L
#define MCI_OPEN_ELEMENT 0x00000200L
#define MCI_OPEN_ALIAS 0x00000400L
#define MCI_OPEN_ELEMENT_ID 0x00000800L
#define MCI_OPEN_TYPE_ID 0x00001000L
#define MCI_OPEN_TYPE 0x00002000L
#define MCI_SEEK_TO_START 0x00000100L
#define MCI_SEEK_TO_END 0x00000200L
#define MCI_STATUS_ITEM 0x00000100L
#define MCI_STATUS_START 0x00000200L
#define MCI_STATUS_LENGTH 0x00000001L
#define MCI_STATUS_POSITION 0x00000002L
#define MCI_STATUS_NUMBER_OF_TRACKS 0x00000003L
#define MCI_STATUS_MODE 0x00000004L
#define MCI_STATUS_MEDIA_PRESENT 0x00000005L
#define MCI_STATUS_TIME_FORMAT 0x00000006L
#define MCI_STATUS_READY 0x00000007L
#define MCI_STATUS_CURRENT_TRACK 0x00000008L
#define MCI_INFO_PRODUCT 0x00000100L
#define MCI_INFO_FILE 0x00000200L
#define MCI_INFO_MEDIA_UPC 0x00000400L
#define MCI_INFO_MEDIA_IDENTITY 0x00000800L
#define MCI_INFO_NAME 0x00001000L
#define MCI_INFO_COPYRIGHT 0x00002000L
#define MCI_GETDEVCAPS_ITEM 0x00000100L
#define MCI_GETDEVCAPS_CAN_RECORD 0x00000001L
#define MCI_GETDEVCAPS_HAS_AUDIO 0x00000002L
#define MCI_GETDEVCAPS_HAS_VIDEO 0x00000003L
#define MCI_GETDEVCAPS_DEVICE_TYPE 0x00000004L
#define MCI_GETDEVCAPS_USES_FILES 0x00000005L
#define MCI_GETDEVCAPS_COMPOUND_DEVICE 0x00000006L
#define MCI_GETDEVCAPS_CAN_EJECT 0x00000007L
#define MCI_GETDEVCAPS_CAN_PLAY 0x00000008L
#define MCI_GETDEVCAPS_CAN_SAVE 0x00000009L
#define MCI_SYSINFO_QUANTITY 0x00000100L
#define MCI_SYSINFO_OPEN 0x00000200L
#define MCI_SYSINFO_NAME 0x00000400L
#define MCI_SYSINFO_INSTALLNAME 0x00000800L
#define MCI_SET_DOOR_OPEN 0x00000100L
#define MCI_SET_DOOR_CLOSED 0x00000200L
#define MCI_SET_TIME_FORMAT 0x00000400L
#define MCI_SET_AUDIO 0x00000800L
#define MCI_SET_VIDEO 0x00001000L
#define MCI_SET_ON 0x00002000L
#define MCI_SET_OFF 0x00004000L
#define MCI_SET_AUDIO_ALL 0x00000000L
#define MCI_SET_AUDIO_LEFT 0x00000001L
#define MCI_SET_AUDIO_RIGHT 0x00000002L
#define MCI_BREAK_KEY 0x00000100L
#define MCI_BREAK_HWND 0x00000200L
#define MCI_BREAK_OFF 0x00000400L
#define MCI_RECORD_INSERT 0x00000100L
#define MCI_RECORD_OVERWRITE 0x00000200L
#define MCI_SAVE_FILE 0x00000100L
#define MCI_LOAD_FILE 0x00000100L
#define MCI_VD_MODE_PARK (MCI_VD_OFFSET + 1)
#define MCI_VD_MEDIA_CLV (MCI_VD_OFFSET + 2)
#define MCI_VD_MEDIA_CAV (MCI_VD_OFFSET + 3)
#define MCI_VD_MEDIA_OTHER (MCI_VD_OFFSET + 4)
#define MCI_VD_FORMAT_TRACK 0x4001
#define MCI_VD_PLAY_REVERSE 0x00010000L
#define MCI_VD_PLAY_FAST 0x00020000L
#define MCI_VD_PLAY_SPEED 0x00040000L
#define MCI_VD_PLAY_SCAN 0x00080000L
#define MCI_VD_PLAY_SLOW 0x00100000L
#define MCI_VD_SEEK_REVERSE 0x00010000L
#define MCI_VD_STATUS_SPEED 0x00004002L
#define MCI_VD_STATUS_FORWARD 0x00004003L
#define MCI_VD_STATUS_MEDIA_TYPE 0x00004004L
#define MCI_VD_STATUS_SIDE 0x00004005L
#define MCI_VD_STATUS_DISC_SIZE 0x00004006L
#define MCI_VD_GETDEVCAPS_CLV 0x00010000L
#define MCI_VD_GETDEVCAPS_CAV 0x00020000L
#define MCI_VD_SPIN_UP 0x00010000L
#define MCI_VD_SPIN_DOWN 0x00020000L
#define MCI_VD_GETDEVCAPS_CAN_REVERSE 0x00004002L
#define MCI_VD_GETDEVCAPS_FAST_RATE 0x00004003L
#define MCI_VD_GETDEVCAPS_SLOW_RATE 0x00004004L
#define MCI_VD_GETDEVCAPS_NORMAL_RATE 0x00004005L
#define MCI_VD_STEP_FRAMES 0x00010000L
#define MCI_VD_STEP_REVERSE 0x00020000L
#define MCI_VD_ESCAPE_STRING 0x00000100L
#define MCI_CDA_STATUS_TYPE_TRACK 0x00004001L
#define MCI_CDA_TRACK_AUDIO (MCI_CD_OFFSET + 0)
#define MCI_CDA_TRACK_OTHER (MCI_CD_OFFSET + 1)
#define MCI_WAVE_PCM (MCI_WAVE_OFFSET + 0)
#define MCI_WAVE_MAPPER (MCI_WAVE_OFFSET + 1)
#define MCI_WAVE_OPEN_BUFFER 0x00010000L
#define MCI_WAVE_SET_FORMATTAG 0x00010000L
#define MCI_WAVE_SET_CHANNELS 0x00020000L
#define MCI_WAVE_SET_SAMPLESPERSEC 0x00040000L
#define MCI_WAVE_SET_AVGBYTESPERSEC 0x00080000L
#define MCI_WAVE_SET_BLOCKALIGN 0x00100000L
#define MCI_WAVE_SET_BITSPERSAMPLE 0x00200000L
#define MCI_WAVE_INPUT 0x00400000L
#define MCI_WAVE_OUTPUT 0x00800000L
#define MCI_WAVE_STATUS_FORMATTAG 0x00004001L
#define MCI_WAVE_STATUS_CHANNELS 0x00004002L
#define MCI_WAVE_STATUS_SAMPLESPERSEC 0x00004003L
#define MCI_WAVE_STATUS_AVGBYTESPERSEC 0x00004004L
#define MCI_WAVE_STATUS_BLOCKALIGN 0x00004005L
#define MCI_WAVE_STATUS_BITSPERSAMPLE 0x00004006L
#define MCI_WAVE_STATUS_LEVEL 0x00004007L
#define MCI_WAVE_SET_ANYINPUT 0x04000000L
#define MCI_WAVE_SET_ANYOUTPUT 0x08000000L
#define MCI_WAVE_GETDEVCAPS_INPUTS 0x00004001L
#define MCI_WAVE_GETDEVCAPS_OUTPUTS 0x00004002L
#define MCI_SEQ_DIV_PPQN (0 + MCI_SEQ_OFFSET)
#define MCI_SEQ_DIV_SMPTE_24 (1 + MCI_SEQ_OFFSET)
#define MCI_SEQ_DIV_SMPTE_25 (2 + MCI_SEQ_OFFSET)
#define MCI_SEQ_DIV_SMPTE_30DROP (3 + MCI_SEQ_OFFSET)
#define MCI_SEQ_DIV_SMPTE_30 (4 + MCI_SEQ_OFFSET)
#define MCI_SEQ_FORMAT_SONGPTR 0x4001
#define MCI_SEQ_FILE 0x4002
#define MCI_SEQ_MIDI 0x4003
#define MCI_SEQ_SMPTE 0x4004
#define MCI_SEQ_NONE 65533
#define MCI_SEQ_MAPPER 65535
#define MCI_SEQ_STATUS_TEMPO 0x00004002L
#define MCI_SEQ_STATUS_PORT 0x00004003L
#define MCI_SEQ_STATUS_SLAVE 0x00004007L
#define MCI_SEQ_STATUS_MASTER 0x00004008L
#define MCI_SEQ_STATUS_OFFSET 0x00004009L
#define MCI_SEQ_STATUS_DIVTYPE 0x0000400AL
#define MCI_SEQ_STATUS_NAME 0x0000400BL
#define MCI_SEQ_STATUS_COPYRIGHT 0x0000400CL
#define MCI_SEQ_SET_TEMPO 0x00010000L
#define MCI_SEQ_SET_PORT 0x00020000L
#define MCI_SEQ_SET_SLAVE 0x00040000L
#define MCI_SEQ_SET_MASTER 0x00080000L
#define MCI_SEQ_SET_OFFSET 0x01000000L
#define MCI_ANIM_OPEN_WS 0x00010000L
#define MCI_ANIM_OPEN_PARENT 0x00020000L
#define MCI_ANIM_OPEN_NOSTATIC 0x00040000L
#define MCI_ANIM_PLAY_SPEED 0x00010000L
#define MCI_ANIM_PLAY_REVERSE 0x00020000L
#define MCI_ANIM_PLAY_FAST 0x00040000L
#define MCI_ANIM_PLAY_SLOW 0x00080000L
#define MCI_ANIM_PLAY_SCAN 0x00100000L
#define MCI_ANIM_STEP_REVERSE 0x00010000L
#define MCI_ANIM_STEP_FRAMES 0x00020000L
#define MCI_ANIM_STATUS_SPEED 0x00004001L
#define MCI_ANIM_STATUS_FORWARD 0x00004002L
#define MCI_ANIM_STATUS_HWND 0x00004003L
#define MCI_ANIM_STATUS_HPAL 0x00004004L
#define MCI_ANIM_STATUS_STRETCH 0x00004005L
#define MCI_ANIM_INFO_TEXT 0x00010000L
#define MCI_ANIM_GETDEVCAPS_CAN_REVERSE 0x00004001L
#define MCI_ANIM_GETDEVCAPS_FAST_RATE 0x00004002L
#define MCI_ANIM_GETDEVCAPS_SLOW_RATE 0x00004003L
#define MCI_ANIM_GETDEVCAPS_NORMAL_RATE 0x00004004L
#define MCI_ANIM_GETDEVCAPS_PALETTES 0x00004006L
#define MCI_ANIM_GETDEVCAPS_CAN_STRETCH 0x00004007L
#define MCI_ANIM_GETDEVCAPS_MAX_WINDOWS 0x00004008L
#define MCI_ANIM_REALIZE_NORM 0x00010000L
#define MCI_ANIM_REALIZE_BKGD 0x00020000L
#define MCI_ANIM_WINDOW_HWND 0x00010000L
#define MCI_ANIM_WINDOW_STATE 0x00040000L
#define MCI_ANIM_WINDOW_TEXT 0x00080000L
#define MCI_ANIM_WINDOW_ENABLE_STRETCH 0x00100000L
#define MCI_ANIM_WINDOW_DISABLE_STRETCH 0x00200000L
#define MCI_ANIM_WINDOW_DEFAULT 0x00000000L
#define MCI_ANIM_RECT 0x00010000L
#define MCI_ANIM_PUT_SOURCE 0x00020000L
#define MCI_ANIM_PUT_DESTINATION 0x00040000L
#define MCI_ANIM_WHERE_SOURCE 0x00020000L
#define MCI_ANIM_WHERE_DESTINATION 0x00040000L
#define MCI_ANIM_UPDATE_HDC 0x00020000L
#define MCI_OVLY_OPEN_WS 0x00010000L
#define MCI_OVLY_OPEN_PARENT 0x00020000L
#define MCI_OVLY_STATUS_HWND 0x00004001L
#define MCI_OVLY_STATUS_STRETCH 0x00004002L
#define MCI_OVLY_INFO_TEXT 0x00010000L
#define MCI_OVLY_GETDEVCAPS_CAN_STRETCH 0x00004001L
#define MCI_OVLY_GETDEVCAPS_CAN_FREEZE 0x00004002L
#define MCI_OVLY_GETDEVCAPS_MAX_WINDOWS 0x00004003L
#define MCI_OVLY_WINDOW_HWND 0x00010000L
#define MCI_OVLY_WINDOW_STATE 0x00040000L
#define MCI_OVLY_WINDOW_TEXT 0x00080000L
#define MCI_OVLY_WINDOW_ENABLE_STRETCH 0x00100000L
#define MCI_OVLY_WINDOW_DISABLE_STRETCH 0x00200000L
#define MCI_OVLY_WINDOW_DEFAULT 0x00000000L
#define MCI_OVLY_RECT 0x00010000L
#define MCI_OVLY_PUT_SOURCE 0x00020000L
#define MCI_OVLY_PUT_DESTINATION 0x00040000L
#define MCI_OVLY_PUT_FRAME 0x00080000L
#define MCI_OVLY_PUT_VIDEO 0x00100000L
#define MCI_OVLY_WHERE_SOURCE 0x00020000L
#define MCI_OVLY_WHERE_DESTINATION 0x00040000L
#define MCI_OVLY_WHERE_FRAME 0x00080000L
#define MCI_OVLY_WHERE_VIDEO 0x00100000L
#define SELECTDIB 41
#define NCBNAMSZ 16
#define MAX_LANA 254
#define NAME_FLAGS_MASK 0x87
#define GROUP_NAME 0x80
#define UNIQUE_NAME 0x00
#define REGISTERING 0x00
#define REGISTERED 0x04
#define DEREGISTERED 0x05
#define DUPLICATE 0x06
#define DUPLICATE_DEREG 0x07
#define LISTEN_OUTSTANDING 0x01
#define CALL_PENDING 0x02
#define SESSION_ESTABLISHED 0x03
#define HANGUP_PENDING 0x04
#define HANGUP_COMPLETE 0x05
#define SESSION_ABORTED 0x06
#define ALL_TRANSPORTS "M\0\0\0"
#define MS_NBF "MNBF"
#define NCBCALL 0x10
#define NCBLISTEN 0x11
#define NCBHANGUP 0x12
#define NCBSEND 0x14
#define NCBRECV 0x15
#define NCBRECVANY 0x16
#define NCBCHAINSEND 0x17
#define NCBDGSEND 0x20
#define NCBDGRECV 0x21
#define NCBDGSENDBC 0x22
#define NCBDGRECVBC 0x23
#define NCBADDNAME 0x30
#define NCBDELNAME 0x31
#define NCBRESET 0x32
#define NCBASTAT 0x33
#define NCBSSTAT 0x34
#define NCBCANCEL 0x35
#define NCBADDGRNAME 0x36
#define NCBENUM 0x37
#define NCBUNLINK 0x70
#define NCBSENDNA 0x71
#define NCBCHAINSENDNA 0x72
#define NCBLANSTALERT 0x73
#define NCBACTION 0x77
#define NCBFINDNAME 0x78
#define NCBTRACE 0x79
#define ASYNCH 0x80
#define NRC_GOODRET 0x00
#define NRC_BUFLEN 0x01
#define NRC_ILLCMD 0x03
#define NRC_CMDTMO 0x05
#define NRC_INCOMP 0x06
#define NRC_BADDR 0x07
#define NRC_SNUMOUT 0x08
#define NRC_NORES 0x09
#define NRC_SCLOSED 0x0a
#define NRC_CMDCAN 0x0b
#define NRC_DUPNAME 0x0d
#define NRC_NAMTFUL 0x0e
#define NRC_ACTSES 0x0f
#define NRC_LOCTFUL 0x11
#define NRC_REMTFUL 0x12
#define NRC_ILLNN 0x13
#define NRC_NOCALL 0x14
#define NRC_NOWILD 0x15
#define NRC_INUSE 0x16
#define NRC_NAMERR 0x17
#define NRC_SABORT 0x18
#define NRC_NAMCONF 0x19
#define NRC_IFBUSY 0x21
#define NRC_TOOMANY 0x22
#define NRC_BRIDGE 0x23
#define NRC_CANOCCR 0x24
#define NRC_CANCEL 0x26
#define NRC_DUPENV 0x30
#define NRC_ENVNOTDEF 0x34
#define NRC_OSRESNOTAV 0x35
#define NRC_MAXAPPS 0x36
#define NRC_NOSAPS 0x37
#define NRC_NORESOURCES 0x38
#define NRC_INVADDRESS 0x39
#define NRC_INVDDID 0x3B
#define NRC_LOCKFAIL 0x3C
#define NRC_OPENERR 0x3f
#define NRC_SYSTEM 0x40
#define NRC_PENDING 0xff
#define IDLFLAG_NONE 0
#define IDLFLAG_FIN 0x1
#define IDLFLAG_FOUT 0x2
#define IDLFLAG_FLCID 0x4
#define IDLFLAG_FRETVAL 0x08
#define DISPATCH_PROPERTYGET 0x2
#define DISPATCH_PROPERTYPUT 0x4
#define DISPATCH_PROPERTYPUTREF 0x8
#define INVOKE_METHOD DISPATCH_METHOD
#define INVOKE_PROPERTYGET DISPATCH_PROPERTYGET
#define INVOKE_PROPERTYPUT DISPATCH_PROPERTYPUT
#define INVOKE_PROPERTYPUTREF DISPATCH_PROPERTYPUTREF
#define FADF_AUTO 0x1
#define FADF_STATIC 0x2
#define FADF_EMBEDDED 0x4
#define FADF_FIXEDSIZE 0x10
#define FADF_RECORD 0x20
#define FADF_HAVEIID 0x40
#define FADF_HAVEVARTYPE 0x80
#define FADF_BSTR 0x100
#define FADF_UNKNOWN 0x200
#define FADF_DISPATCH 0x400
#define FADF_VARIANT 0x800
#define FADF_RESERVED 0xf0e8
#define VARFLAG_FREADONLY 1
#define VARFLAG_FSOURCE 0x2
#define VARFLAG_FBINDABLE 0x4
#define VARFLAG_FREQUESTEDIT 0x8
#define VARFLAG_FDISPLAYBIND 0x10
#define VARFLAG_FDEFAULTBIND 0x20
#define VARFLAG_FHIDDEN 0x40
#define VARFLAG_FRESTRICTED 0x80
#define VARFLAG_FDEFAULTCOLLELEM 0x100
#define VARFLAG_FUIDEFAULT 0x200
#define VARFLAG_FNONBROWSABLE 0x400
#define VARFLAG_FREPLACEABLE 0x800
#define VARFLAG_FIMMEDIATEBIND 0x1000
#define TYPEFLAG_FAPPOBJECT 0x1
#define TYPEFLAG_FCANCREATE 0x2
#define TYPEFLAG_FLICENSED 0x4
#define TYPEFLAG_FPREDECLID 0x8
#define TYPEFLAG_FHIDDEN 0x10
#define TYPEFLAG_FCONTROL 0x20
#define TYPEFLAG_FDUAL 0x40
#define TYPEFLAG_FNONEXTENSIBLE 0x80
#define TYPEFLAG_FOLEAUTOMATION 0x100
#define TYPEFLAG_FRESTRICTED 0x200
#define TYPEFLAG_FAGGREGATABLE 0x400
#define TYPEFLAG_FREPLACEABLE 0x800
#define TYPEFLAG_FDISPATCHABLE 0x1000
#define TYPEFLAG_FREVERSEBIND 0x2000
#define TYPEFLAG_FPROXY 0x4000
#define FUNCFLAG_FRESTRICTED 0x1
#define FUNCFLAG_FSOURCE 0x2
#define FUNCFLAG_FBINDABLE 0x4
#define FUNCFLAG_FREQUESTEDIT 0x8
#define FUNCFLAG_FDISPLAYBIND 0x10
#define FUNCFLAG_FDEFAULTBIND 0x20
#define FUNCFLAG_FHIDDEN 0x40
#define FUNCFLAG_FUSESGETLASTERROR 0x80
#define FUNCFLAG_FDEFAULTCOLLELEM 0x100
#define FUNCFLAG_FUIDEFAULT 0x200
#define FUNCFLAG_FNONBROWSABLE 0x400
#define FUNCFLAG_FREPLACEABLE 0x800
#define FUNCFLAG_FIMMEDIATEBIND 0x1000
#define VT_EMPTY 0
#define VT_NULL 1
#define VT_I2 2
#define VT_I4 3
#define VT_R4 4
#define VT_R8 5
#define VT_CY 6
#define VT_DATE 7
#define VT_BSTR 8
#define VT_DISPATCH 9
#define VT_ERROR 10
#define VT_BOOL 11
#define VT_VARIANT 12
#define VT_UNKNOWN 13
#define VT_DECIMAL 14
#define VT_I1 16
#define VT_UI1 17
#define VT_UI2 18
#define VT_UI4 19
#define VT_I8 20
#define VT_UI8 21
#define VT_INT 22
#define VT_UINT 23
#define VT_VOID 24
#define VT_HRESULT 25
#define VT_PTR 26
#define VT_SAFEARRAY 27
#define VT_CARRAY 28
#define VT_USERDEFINED 29
#define VT_LPSTR 30
#define VT_LPWSTR 31
#define VT_RECORD 36
#define VT_INT_PTR 37
#define VT_UINT_PTR 38
#define VT_FILETIME 64
#define VT_BLOB 65
#define VT_STREAM 66
#define VT_STORAGE 67
#define VT_STREAMED_OBJECT 68
#define VT_STORED_OBJECT 69
#define VT_BLOB_OBJECT 70
#define VT_CF 71
#define VT_CLSID 72
#define VT_VERSIONED_STREAM 73
#define VT_VECTOR 0x1000
#define VT_ARRAY 0x2000
#define VT_BYREF 0x4000
#define VT_RESERVED 0x8000
#define VT_ILLEGAL 0xFFFF
#define VT_ILLEGALMASKED 0xFFF
#define VT_TYPEMASK 0xFFF
#define DISPID_VALUE ( 0 )
#define DISPID_PROPERTYPUT ( -3 )
#define DISPID_NEWENUM ( -4 )
#define DISPID_EVALUATE ( -5 )
#define DISPID_CONSTRUCTOR ( -6 )
#define DISPID_DESTRUCTOR ( -7 )
#define DISPID_COLLECT ( -8 )
#define STDOLE_MAJORVERNUM 0x1
#define STDOLE_MINORVERNUM 0x0
#define STDOLE_LCID 0x0000
#define VARIANT_NOVALUEPROP 1
#define VARIANT_ALPHABOOL 0x02
#define VARIANT_NOUSEROVERRIDE 0x04
#define VAR_TIMEVALUEONLY 0x0001
#define VAR_DATEVALUEONLY 0x0002
#define ID_DEFAULTINST -2
#define ACTIVEOBJECT_STRONG 0x0
#define ACTIVEOBJECT_WEAK 0x1
#define triUnchecked 0
#define triChecked 1
#define triGray 2
#define VT_STREAMED_PROPSET 73
#define VT_STORED_PROPSET 74
#define VT_BLOB_PROPSET 75
#define VT_VERBOSE_ENUM 76
#define VT_COLOR 3
#define VT_XPOS_PIXELS 3
#define VT_YPOS_PIXELS 3
#define VT_XSIZE_PIXELS 3
#define VT_YSIZE_PIXELS 3
#define VT_XPOS_HIMETRIC 3
#define VT_YPOS_HIMETRIC 3
#define VT_XSIZE_HIMETRIC 3
#define VT_YSIZE_HIMETRIC 3
#define VT_TRISTATE 2
#define VT_OPTEXCLUSIVE 11
#define VT_FONT 9
#define VT_PICTURE 9
#define VT_HANDLE 3
#define OCM__BASE (WM_USER+0x1c00)
#define WM_COMMAND 0x0111
#define OCM_COMMAND (OCM__BASE + WM_COMMAND)
#define WM_CTLCOLORBTN 0x0135
#define OCM_CTLCOLORBTN (OCM__BASE + WM_CTLCOLORBTN)
#define WM_CTLCOLOREDIT 0x0133
#define OCM_CTLCOLOREDIT (OCM__BASE + WM_CTLCOLOREDIT)
#define WM_CTLCOLORDLG 0x0136
#define OCM_CTLCOLORDLG (OCM__BASE + WM_CTLCOLORDLG)
#define WM_CTLCOLORLISTBOX 0x0134
#define OCM_CTLCOLORLISTBOX (OCM__BASE + WM_CTLCOLORLISTBOX)
#define WM_CTLCOLORMSGBOX 0x0132
#define OCM_CTLCOLORMSGBOX (OCM__BASE + WM_CTLCOLORMSGBOX)
#define WM_CTLCOLORSCROLLBAR 0x0137
#define OCM_CTLCOLORSCROLLBAR (OCM__BASE + WM_CTLCOLORSCROLLBAR)
#define WM_CTLCOLORSTATIC 0x0138
#define OCM_CTLCOLORSTATIC (OCM__BASE + WM_CTLCOLORSTATIC)
#define WM_DRAWITEM 0x002B
#define OCM_DRAWITEM (OCM__BASE + WM_DRAWITEM)
#define WM_MEASUREITEM 0x002C
#define OCM_MEASUREITEM (OCM__BASE + WM_MEASUREITEM)
#define WM_DELETEITEM 0x002D
#define OCM_DELETEITEM (OCM__BASE + WM_DELETEITEM)
#define WM_VKEYTOITEM 0x002E
#define OCM_VKEYTOITEM (OCM__BASE + WM_VKEYTOITEM)
#define WM_CHARTOITEM 0x002F
#define OCM_CHARTOITEM (OCM__BASE + WM_CHARTOITEM)
#define WM_COMPAREITEM 0x0039
#define OCM_COMPAREITEM (OCM__BASE + WM_COMPAREITEM)
#define WM_HSCROLL 0x0114
#define OCM_HSCROLL (OCM__BASE + WM_HSCROLL)
#define WM_VSCROLL 0x0115
#define OCM_VSCROLL (OCM__BASE + WM_VSCROLL)
#define WM_PARENTNOTIFY 0x0210
#define OCM_PARENTNOTIFY (OCM__BASE + WM_PARENTNOTIFY)
#define CTRLINFO_EATS_RETURN 1
#define CTRLINFO_EATS_ESCAPE 2
#define XFORMCOORDS_POSITION 0x1
#define XFORMCOORDS_SIZE 0x2
#define XFORMCOORDS_HIMETRICTOCONTAINER 0x4
#define XFORMCOORDS_CONTAINERTOHIMETRIC 0x8
#define PROPPAGESTATUS_DIRTY 0x1
#define PROPPAGESTATUS_VALIDATE 0x2
#define PICTURE_SCALABLE 0x1l
#define PICTURE_TRANSPARENT 0x2l
#define PICTYPE_UNINITIALIZED DWORD(_cast, 0xffffffff)
#define PICTYPE_NONE 0
#define PICTYPE_BITMAP 1
#define PICTYPE_METAFILE 2
#define PICTYPE_ICON 3
#define DISPID_AUTOSIZE (-500)
#define DISPID_BACKCOLOR (-501)
#define DISPID_BACKSTYLE (-502)
#define DISPID_BORDERCOLOR (-503)
#define DISPID_BORDERSTYLE (-504)
#define DISPID_BORDERWIDTH (-505)
#define DISPID_DRAWMODE (-507)
#define DISPID_DRAWSTYLE (-508)
#define DISPID_DRAWWIDTH (-509)
#define DISPID_FILLCOLOR (-510)
#define DISPID_FILLSTYLE (-511)
#define DISPID_FONT (-512)
#define DISPID_FORECOLOR (-513)
#define DISPID_ENABLED (-514)
#define DISPID_HWND (-515)
#define DISPID_TABSTOP (-516)
#define DISPID_TEXT (-517)
#define DISPID_CAPTION (-518)
#define DISPID_BORDERVISIBLE (-519)
#define DISPID_REFRESH (-550)
#define DISPID_DOCLICK (-551)
#define DISPID_ABOUTBOX (-552)
#define DISPID_CLICK (-600)
#define DISPID_DBLCLICK (-601)
#define DISPID_KEYDOWN (-602)
#define DISPID_KEYPRESS (-603)
#define DISPID_KEYUP (-604)
#define DISPID_MOUSEDOWN (-605)
#define DISPID_MOUSEMOVE (-606)
#define DISPID_MOUSEUP (-607)
#define DISPID_ERROREVENT (-608)
#define DISPID_AMBIENT_BACKCOLOR (-701)
#define DISPID_AMBIENT_DISPLAYNAME (-702)
#define DISPID_AMBIENT_FONT (-703)
#define DISPID_AMBIENT_FORECOLOR (-704)
#define DISPID_AMBIENT_LOCALEID (-705)
#define DISPID_AMBIENT_MESSAGEREFLECT (-706)
#define DISPID_AMBIENT_SCALEUNITS (-707)
#define DISPID_AMBIENT_TEXTALIGN (-708)
#define DISPID_AMBIENT_USERMODE (-709)
#define DISPID_AMBIENT_UIDEAD (-710)
#define DISPID_AMBIENT_SHOWGRABHANDLES (-711)
#define DISPID_AMBIENT_SHOWHATCHING (-712)
#define DISPID_AMBIENT_DISPLAYASDEFAULT (-713)
#define DISPID_AMBIENT_SUPPORTSMNEMONICS (-714)
#define DISPID_AMBIENT_AUTOCLIP (-715)
#define DISPID_FONT_NAME 0
#define DISPID_FONT_SIZE 2
#define DISPID_FONT_BOLD 3
#define DISPID_FONT_ITALIC 4
#define DISPID_FONT_UNDER 5
#define DISPID_FONT_STRIKE 6
#define DISPID_FONT_WEIGHT 7
#define DISPID_FONT_CHARSET 8
#define DISPID_PICT_HANDLE 0
#define DISPID_PICT_HPAL 2
#define DISPID_PICT_TYPE 3
#define DISPID_PICT_WIDTH 4
#define DISPID_PICT_HEIGHT 5
#define DISPID_PICT_RENDER 6
#define STDOLE_TLB "stdole32.tlb"
#define STDTYPE_TLB "oc30d.dll"
#define LPD_DOUBLEBUFFER 0x00000001
#define LPD_STEREO 0x00000002
#define LPD_SUPPORT_GDI 0x00000010
#define LPD_SUPPORT_OPENGL 0x00000020
#define LPD_SHARE_DEPTH 0x00000040
#define LPD_SHARE_STENCIL 0x00000080
#define LPD_SHARE_ACCUM 0x00000100
#define LPD_SWAP_EXCHANGE 0x00000200
#define LPD_SWAP_COPY 0x00000400
#define LPD_TRANSPARENT 0x00001000
#define LPD_TYPE_RGBA 0
#define LPD_TYPE_COLORINDEX 1
#define WGL_SWAP_MAIN_PLANE 0x00000001
#define WGL_SWAP_OVERLAY1 0x00000002
#define WGL_SWAP_OVERLAY2 0x00000004
#define WGL_SWAP_OVERLAY3 0x00000008
#define WGL_SWAP_OVERLAY4 0x00000010
#define WGL_SWAP_OVERLAY5 0x00000020
#define WGL_SWAP_OVERLAY6 0x00000040
#define WGL_SWAP_OVERLAY7 0x00000080
#define WGL_SWAP_OVERLAY8 0x00000100
#define WGL_SWAP_OVERLAY9 0x00000200
#define WGL_SWAP_OVERLAY10 0x00000400
#define WGL_SWAP_OVERLAY11 0x00000800
#define WGL_SWAP_OVERLAY12 0x00001000
#define WGL_SWAP_OVERLAY13 0x00002000
#define WGL_SWAP_OVERLAY14 0x00004000
#define WGL_SWAP_OVERLAY15 0x00008000
#define WGL_SWAP_UNDERLAY1 0x00010000
#define WGL_SWAP_UNDERLAY2 0x00020000
#define WGL_SWAP_UNDERLAY3 0x00040000
#define WGL_SWAP_UNDERLAY4 0x00080000
#define WGL_SWAP_UNDERLAY5 0x00100000
#define WGL_SWAP_UNDERLAY6 0x00200000
#define WGL_SWAP_UNDERLAY7 0x00400000
#define WGL_SWAP_UNDERLAY8 0x00800000
#define WGL_SWAP_UNDERLAY9 0x01000000
#define WGL_SWAP_UNDERLAY10 0x02000000
#define WGL_SWAP_UNDERLAY11 0x04000000
#define WGL_SWAP_UNDERLAY12 0x08000000
#define WGL_SWAP_UNDERLAY13 0x10000000
#define WGL_SWAP_UNDERLAY14 0x20000000
#define WGL_SWAP_UNDERLAY15 0x40000000
#define RAS_MaxDeviceType 16
#define RAS_MaxPhoneNumber 128
#define RAS_MaxIpAddress 15
#define RAS_MaxIpxAddress 21
#define RAS_MaxEntryName 256
#define RAS_MaxDeviceName 128
#define RAS_MaxCallbackNumber RAS_MaxPhoneNumber
#define RAS_MaxAreaCode 10
#define RAS_MaxPadType 32
#define RAS_MaxX25Address 200
#define RAS_MaxFacilities 200
#define RAS_MaxUserData 200
#define RAS_MaxReplyMessage 1024
#define RAS_MaxDnsSuffix 256
#define RASCF_AllUsers 0x00000001
#define RASCF_GlobalCreds 0x00000002
#define RASCS_PAUSED 0x1000
#define RASCS_DONE 0x2000
#define RASCS_OpenPort 0
#define RASCS_PortOpened 1
#define RASCS_ConnectDevice 2
#define RASCS_DeviceConnected 3
#define RASCS_AllDevicesConnected 4
#define RASCS_Authenticate 5
#define RASCS_AuthNotify 6
#define RASCS_AuthRetry 7
#define RASCS_AuthCallback 8
#define RASCS_AuthChangePassword 9
#define RASCS_AuthProject 10
#define RASCS_AuthLinkSpeed 11
#define RASCS_AuthAck 12
#define RASCS_ReAuthenticate 13
#define RASCS_Authenticated 14
#define RASCS_PrepareForCallback 15
#define RASCS_WaitForModemReset 16
#define RASCS_WaitForCallback 17
#define RASCS_Projected 18
#define RASCS_StartAuthentication 19
#define RASCS_CallbackComplete 20
#define RASCS_LogonNetwork 21
#define RASCS_SubEntryConnected 22
#define RASCS_SubEntryDisconnected 23
#define RASCS_Interactive RASCS_PAUSED
#define RASCS_RetryAuthentication 24
#define RASCS_CallbackSetByCaller 25
#define RASCS_PasswordExpired 26
#define RASCS_InvokeEapUI 27
#define RASCS_Connected RASCS_DONE
#define RASCS_Disconnected RASCS_DONE+1
#define RDEOPT_UsePrefixSuffix 0x00000001
#define RDEOPT_PausedStates 0x00000002
#define RDEOPT_IgnoreModemSpeaker 0x00000004
#define RDEOPT_SetModemSpeaker 0x00000008
#define RDEOPT_IgnoreSoftwareCompression 0x00000010
#define RDEOPT_SetSoftwareCompression 0x00000020
#define RDEOPT_DisableConnectedUI 0x00000040
#define RDEOPT_DisableReconnectUI 0x00000080
#define RDEOPT_DisableReconnect 0x00000100
#define RDEOPT_NoUser 0x00000200
#define RDEOPT_PauseOnScript 0x00000400
#define RDEOPT_Router 0x00000800
#define RDEOPT_CustomDial 0x00001000
#define RDEOPT_UseCustomScripting 0x00002000
#define REN_User 0x00000000
#define REN_AllUsers 0x00000001
#define RASP_Amb 0x10000
#define RASP_PppNbf 0x803F
#define RASP_PppIpx 0x802B
#define RASP_PppIp 0x8021
#define RASP_PppCcp 0x80FD
#define RASP_PppLcp 0xC021
#define RASP_Slip 0x20000
#define RASLCPAP_PAP 0xC023
#define RASLCPAP_SPAP 0xC027
#define RASLCPAP_CHAP 0xC223
#define RASLCPAP_EAP 0xC227
#define RASLCPAD_CHAP_MD5 0x05
#define RASLCPAD_CHAP_MS 0x80
#define RASLCPAD_CHAP_MSV2 0x81
#define RASLCPO_PFC 0x00000001
#define RASLCPO_ACFC 0x00000002
#define RASLCPO_SSHF 0x00000004
#define RASLCPO_DES_56 0x00000008
#define RASLCPO_3_DES 0x00000010
#define RASDIALEVENT "RasDialEvent"
#define WM_RASDIALEVENT 0xCCCD
#define ET_None 0
#define ET_Require 1
#define ET_RequireMax 2
#define ET_Optional 3
#define VS_Default 0
#define VS_PptpOnly 1
#define VS_PptpFirst 2
#define VS_L2tpOnly 3
#define VS_L2tpFirst 4
#define RASEO_UseCountryAndAreaCodes 0x00000001
#define RASEO_SpecificIpAddr 0x00000002
#define RASEO_SpecificNameServers 0x00000004
#define RASEO_IpHeaderCompression 0x00000008
#define RASEO_RemoteDefaultGateway 0x00000010
#define RASEO_DisableLcpExtensions 0x00000020
#define RASEO_TerminalBeforeDial 0x00000040
#define RASEO_TerminalAfterDial 0x00000080
#define RASEO_ModemLights 0x00000100
#define RASEO_SwCompression 0x00000200
#define RASEO_RequireEncryptedPw 0x00000400
#define RASEO_RequireMsEncryptedPw 0x00000800
#define RASEO_RequireDataEncryption 0x00001000
#define RASEO_NetworkLogon 0x00002000
#define RASEO_UseLogonCredentials 0x00004000
#define RASEO_PromoteAlternates 0x00008000
#define RASEO_SecureLocalFiles 0x00010000
#define RASEO_RequireEAP 0x00020000
#define RASEO_RequirePAP 0x00040000
#define RASEO_RequireSPAP 0x00080000
#define RASEO_Custom 0x00100000
#define RASEO_PreviewPhoneNumber 0x00200000
#define RASEO_SharedPhoneNumbers 0x00800000
#define RASEO_PreviewUserPw 0x01000000
#define RASEO_PreviewDomain 0x02000000
#define RASEO_ShowDialingProgress 0x04000000
#define RASEO_RequireCHAP 0x08000000
#define RASEO_RequireMsCHAP 0x10000000
#define RASEO_RequireMsCHAP2 0x20000000
#define RASEO_RequireW95MSCHAP 0x40000000
#define RASEO_CustomScript 0x80000000
#define RASEO2_SecureFileAndPrint 0x00000001
#define RASEO2_SecureClientForMSNet 0x00000002
#define RASEO2_DontNegotiateMultilink 0x00000004
#define RASEO2_DontUseRasCredentials 0x00000008
#define RASEO2_UsePreSharedKey 0x00000010
#define RASEO2_Internet 0x00000020
#define RASEO2_DisableNbtOverIP 0x00000040
#define RASEO2_UseGlobalDeviceSettings 0x00000080
#define RASEO2_ReconnectIfDropped 0x00000100
#define RASEO2_SharePhoneNumbers 0x00000200
#define RASNP_NetBEUI 0x00000001
#define RASNP_Ipx 0x00000002
#define RASNP_Ip 0x00000004
#define RASFP_Ppp 0x00000001
#define RASFP_Slip 0x00000002
#define RASFP_Ras 0x00000004
#define RASDT_Modem "modem"
#define RASDT_Isdn "isdn"
#define RASDT_X25 "x25"
#define RASDT_Vpn "vpn"
#define RASDT_Pad "pad"
#define RASDT_Generic "GENERIC"
#define RASDT_Serial "SERIAL"
#define RASDT_FrameRelay "FRAMERELAY"
#define RASDT_Atm "ATM"
#define RASDT_Sonet "SONET"
#define RASDT_SW56 "SW56"
#define RASDT_Irda "IRDA"
#define RASDT_Parallel "PARALLEL"
#define RASDT_PPPoE "PPPoE"
#define RASET_Phone 1
#define RASET_Vpn 2
#define RASET_Direct 3
#define RASET_Internet 4
#define RASET_Broadband 5
#define RASCN_Connection 0x00000001
#define RASCN_Disconnection 0x00000002
#define RASCN_BandwidthAdded 0x00000004
#define RASCN_BandwidthRemoved 0x00000008
#define RASEDM_DialAll 1
#define RASEDM_DialAsNeeded 2
#define RASIDS_Disabled 0xffffffff
#define RASIDS_UseGlobalValue 0
#define RASADFLG_PositionDlg 0x00000001
#define RASCM_UserName 0x00000001
#define RASCM_Password 0x00000002
#define RASCM_Domain 0x00000004
#define RASCM_DefaultCreds 0x00000008
#define RASCM_PreSharedKey 0x00000010
#define RASCM_ServerPreSharedKey 0x00000020
#define RASCM_DDMPreSharedKey 0x00000040
#define RASADP_DisableConnectionQuery 0
#define RASADP_LoginSessionDisable 1
#define RASADP_SavedAddressesLimit 2
#define RASADP_FailedConnectionTimeout 3
#define RASADP_ConnectionQueryTimeout 4
#define RASEAPF_NonInteractive 0x00000002
#define RASEAPF_Logon 0x00000004
#define RASEAPF_Preview 0x00000008
#define RASBASE 600
#define SUCCESS 0
#define PENDING (RASBASE+0)
#define ERROR_INVALID_PORT_HANDLE (RASBASE+1)
#define ERROR_PORT_ALREADY_OPEN (RASBASE+2)
#define ERROR_BUFFER_TOO_SMALL (RASBASE+3)
#define ERROR_WRONG_INFO_SPECIFIED (RASBASE+4)
#define ERROR_CANNOT_SET_PORT_INFO (RASBASE+5)
#define ERROR_PORT_NOT_CONNECTED (RASBASE+6)
#define ERROR_EVENT_INVALID (RASBASE+7)
#define ERROR_DEVICE_DOES_NOT_EXIST (RASBASE+8)
#define ERROR_DEVICETYPE_DOES_NOT_EXIST (RASBASE+9)
#define ERROR_BUFFER_INVALID (RASBASE+10)
#define ERROR_ROUTE_NOT_AVAILABLE (RASBASE+11)
#define ERROR_ROUTE_NOT_ALLOCATED (RASBASE+12)
#define ERROR_INVALID_COMPRESSION_SPECIFIED (RASBASE+13)
#define ERROR_OUT_OF_BUFFERS (RASBASE+14)
#define ERROR_PORT_NOT_FOUND (RASBASE+15)
#define ERROR_ASYNC_REQUEST_PENDING (RASBASE+16)
#define ERROR_ALREADY_DISCONNECTING (RASBASE+17)
#define ERROR_PORT_NOT_OPEN (RASBASE+18)
#define ERROR_PORT_DISCONNECTED (RASBASE+19)
#define ERROR_NO_ENDPOINTS (RASBASE+20)
#define ERROR_CANNOT_OPEN_PHONEBOOK (RASBASE+21)
#define ERROR_CANNOT_LOAD_PHONEBOOK (RASBASE+22)
#define ERROR_CANNOT_FIND_PHONEBOOK_ENTRY (RASBASE+23)
#define ERROR_CANNOT_WRITE_PHONEBOOK (RASBASE+24)
#define ERROR_CORRUPT_PHONEBOOK (RASBASE+25)
#define ERROR_CANNOT_LOAD_STRING (RASBASE+26)
#define ERROR_KEY_NOT_FOUND (RASBASE+27)
#define ERROR_DISCONNECTION (RASBASE+28)
#define ERROR_REMOTE_DISCONNECTION (RASBASE+29)
#define ERROR_HARDWARE_FAILURE (RASBASE+30)
#define ERROR_USER_DISCONNECTION (RASBASE+31)
#define ERROR_INVALID_SIZE (RASBASE+32)
#define ERROR_PORT_NOT_AVAILABLE (RASBASE+33)
#define ERROR_CANNOT_PROJECT_CLIENT (RASBASE+34)
#define ERROR_UNKNOWN (RASBASE+35)
#define ERROR_WRONG_DEVICE_ATTACHED (RASBASE+36)
#define ERROR_BAD_STRING (RASBASE+37)
#define ERROR_REQUEST_TIMEOUT (RASBASE+38)
#define ERROR_CANNOT_GET_LANA (RASBASE+39)
#define ERROR_NETBIOS_ERROR (RASBASE+40)
#define ERROR_SERVER_OUT_OF_RESOURCES (RASBASE+41)
#define ERROR_NAME_EXISTS_ON_NET (RASBASE+42)
#define ERROR_SERVER_GENERAL_NET_FAILURE (RASBASE+43)
#define WARNING_MSG_ALIAS_NOT_ADDED (RASBASE+44)
#define ERROR_AUTH_INTERNAL (RASBASE+45)
#define ERROR_RESTRICTED_LOGON_HOURS (RASBASE+46)
#define ERROR_ACCT_DISABLED (RASBASE+47)
#define ERROR_PASSWD_EXPIRED (RASBASE+48)
#define ERROR_NO_DIALIN_PERMISSION (RASBASE+49)
#define ERROR_SERVER_NOT_RESPONDING (RASBASE+50)
#define ERROR_FROM_DEVICE (RASBASE+51)
#define ERROR_UNRECOGNIZED_RESPONSE (RASBASE+52)
#define ERROR_MACRO_NOT_FOUND (RASBASE+53)
#define ERROR_MACRO_NOT_DEFINED (RASBASE+54)
#define ERROR_MESSAGE_MACRO_NOT_FOUND (RASBASE+55)
#define ERROR_DEFAULTOFF_MACRO_NOT_FOUND (RASBASE+56)
#define ERROR_FILE_COULD_NOT_BE_OPENED (RASBASE+57)
#define ERROR_DEVICENAME_TOO_LONG (RASBASE+58)
#define ERROR_DEVICENAME_NOT_FOUND (RASBASE+59)
#define ERROR_NO_RESPONSES (RASBASE+60)
#define ERROR_NO_COMMAND_FOUND (RASBASE+61)
#define ERROR_WRONG_KEY_SPECIFIED (RASBASE+62)
#define ERROR_UNKNOWN_DEVICE_TYPE (RASBASE+63)
#define ERROR_ALLOCATING_MEMORY (RASBASE+64)
#define ERROR_PORT_NOT_CONFIGURED (RASBASE+65)
#define ERROR_DEVICE_NOT_READY (RASBASE+66)
#define ERROR_READING_INI_FILE (RASBASE+67)
#define ERROR_NO_CONNECTION (RASBASE+68)
#define ERROR_BAD_USAGE_IN_INI_FILE (RASBASE+69)
#define ERROR_READING_SECTIONNAME (RASBASE+70)
#define ERROR_READING_DEVICETYPE (RASBASE+71)
#define ERROR_READING_DEVICENAME (RASBASE+72)
#define ERROR_READING_USAGE (RASBASE+73)
#define ERROR_READING_MAXCONNECTBPS (RASBASE+74)
#define ERROR_READING_MAXCARRIERBPS (RASBASE+75)
#define ERROR_LINE_BUSY (RASBASE+76)
#define ERROR_VOICE_ANSWER (RASBASE+77)
#define ERROR_NO_ANSWER (RASBASE+78)
#define ERROR_NO_CARRIER (RASBASE+79)
#define ERROR_NO_DIALTONE (RASBASE+80)
#define ERROR_IN_COMMAND (RASBASE+81)
#define ERROR_WRITING_SECTIONNAME (RASBASE+82)
#define ERROR_WRITING_DEVICETYPE (RASBASE+83)
#define ERROR_WRITING_DEVICENAME (RASBASE+84)
#define ERROR_WRITING_MAXCONNECTBPS (RASBASE+85)
#define ERROR_WRITING_MAXCARRIERBPS (RASBASE+86)
#define ERROR_WRITING_USAGE (RASBASE+87)
#define ERROR_WRITING_DEFAULTOFF (RASBASE+88)
#define ERROR_READING_DEFAULTOFF (RASBASE+89)
#define ERROR_EMPTY_INI_FILE (RASBASE+90)
#define ERROR_AUTHENTICATION_FAILURE (RASBASE+91)
#define ERROR_PORT_OR_DEVICE (RASBASE+92)
#define ERROR_NOT_BINARY_MACRO (RASBASE+93)
#define ERROR_DCB_NOT_FOUND (RASBASE+94)
#define ERROR_STATE_MACHINES_NOT_STARTED (RASBASE+95)
#define ERROR_STATE_MACHINES_ALREADY_STARTED (RASBASE+96)
#define ERROR_PARTIAL_RESPONSE_LOOPING (RASBASE+97)
#define ERROR_UNKNOWN_RESPONSE_KEY (RASBASE+98)
#define ERROR_RECV_BUF_FULL (RASBASE+99)
#define ERROR_CMD_TOO_LONG (RASBASE+100)
#define ERROR_UNSUPPORTED_BPS (RASBASE+101)
#define ERROR_UNEXPECTED_RESPONSE (RASBASE+102)
#define ERROR_INTERACTIVE_MODE (RASBASE+103)
#define ERROR_BAD_CALLBACK_NUMBER (RASBASE+104)
#define ERROR_INVALID_AUTH_STATE (RASBASE+105)
#define ERROR_WRITING_INITBPS (RASBASE+106)
#define ERROR_X25_DIAGNOSTIC (RASBASE+107)
#define ERROR_ACCT_EXPIRED (RASBASE+108)
#define ERROR_CHANGING_PASSWORD (RASBASE+109)
#define ERROR_OVERRUN (RASBASE+110)
#define ERROR_RASMAN_CANNOT_INITIALIZE (RASBASE+111)
#define ERROR_BIPLEX_PORT_NOT_AVAILABLE (RASBASE+112)
#define ERROR_NO_ACTIVE_ISDN_LINES (RASBASE+113)
#define ERROR_NO_ISDN_CHANNELS_AVAILABLE (RASBASE+114)
#define ERROR_TOO_MANY_LINE_ERRORS (RASBASE+115)
#define ERROR_IP_CONFIGURATION (RASBASE+116)
#define ERROR_NO_IP_ADDRESSES (RASBASE+117)
#define ERROR_PPP_TIMEOUT (RASBASE+118)
#define ERROR_PPP_REMOTE_TERMINATED (RASBASE+119)
#define ERROR_PPP_NO_PROTOCOLS_CONFIGURED (RASBASE+120)
#define ERROR_PPP_NO_RESPONSE (RASBASE+121)
#define ERROR_PPP_INVALID_PACKET (RASBASE+122)
#define ERROR_PHONE_NUMBER_TOO_LONG (RASBASE+123)
#define ERROR_IPXCP_NO_DIALOUT_CONFIGURED (RASBASE+124)
#define ERROR_IPXCP_NO_DIALIN_CONFIGURED (RASBASE+125)
#define ERROR_IPXCP_DIALOUT_ALREADY_ACTIVE (RASBASE+126)
#define ERROR_ACCESSING_TCPCFGDLL (RASBASE+127)
#define ERROR_NO_IP_RAS_ADAPTER (RASBASE+128)
#define ERROR_SLIP_REQUIRES_IP (RASBASE+129)
#define ERROR_PROJECTION_NOT_COMPLETE (RASBASE+130)
#define ERROR_PROTOCOL_NOT_CONFIGURED (RASBASE+131)
#define ERROR_PPP_NOT_CONVERGING (RASBASE+132)
#define ERROR_PPP_CP_REJECTED (RASBASE+133)
#define ERROR_PPP_LCP_TERMINATED (RASBASE+134)
#define ERROR_PPP_REQUIRED_ADDRESS_REJECTED (RASBASE+135)
#define ERROR_PPP_NCP_TERMINATED (RASBASE+136)
#define ERROR_PPP_LOOPBACK_DETECTED (RASBASE+137)
#define ERROR_PPP_NO_ADDRESS_ASSIGNED (RASBASE+138)
#define ERROR_CANNOT_USE_LOGON_CREDENTIALS (RASBASE+139)
#define ERROR_TAPI_CONFIGURATION (RASBASE+140)
#define ERROR_NO_LOCAL_ENCRYPTION (RASBASE+141)
#define ERROR_NO_REMOTE_ENCRYPTION (RASBASE+142)
#define ERROR_REMOTE_REQUIRES_ENCRYPTION (RASBASE+143)
#define ERROR_IPXCP_NET_NUMBER_CONFLICT (RASBASE+144)
#define ERROR_INVALID_SMM (RASBASE+145)
#define ERROR_SMM_UNINITIALIZED (RASBASE+146)
#define ERROR_NO_MAC_FOR_PORT (RASBASE+147)
#define ERROR_SMM_TIMEOUT (RASBASE+148)
#define ERROR_BAD_PHONE_NUMBER (RASBASE+149)
#define ERROR_WRONG_MODULE (RASBASE+150)
#define ERROR_INVALID_CALLBACK_NUMBER (RASBASE+151)
#define RASBASEEND (RASBASE+151)
#define SECURITYMSG_SUCCESS 1
#define SECURITYMSG_FAILURE 2
#define SECURITYMSG_ERROR 3
#define RASPBDEVENT_AddEntry 1
#define RASPBDEVENT_EditEntry 2
#define RASPBDEVENT_RemoveEntry 3
#define RASPBDEVENT_DialEntry 4
#define RASPBDEVENT_EditGlobals 5
#define RASPBDEVENT_NoUser 6
#define RASPBDEVENT_NoUserEdit 7
#define RASPBDFLAG_PositionDlg 0x00000001
#define RASPBDFLAG_ForceCloseOnDial 0x00000002
#define RASPBDFLAG_NoUser 0x00000010
#define RASPBDFLAG_UpdateDefaults 0x80000000
#define RASEDFLAG_PositionDlg 0x00000001
#define RASEDFLAG_NewEntry 0x00000002
#define RASEDFLAG_CloneEntry 0x00000004
#define RASEDFLAG_NoRename 0x00000008
#define RASDDFLAG_PositionDlg 0x00000001
#define RASMDPAGE_Status 0
#define RASMDPAGE_Summary 1
#define RASMDPAGE_Preferences 2
#define RASMDFLAG_PositionDlg 0x00000001
#define RASMDFLAG_UpdateDefaults 0x80000000
#define RASSAPI_MAX_PHONENUMBER_SIZE 128
#define RASSAPI_MAX_MEDIA_NAME 16
#define RASSAPI_MAX_PORT_NAME 16
#define RASSAPI_MAX_DEVICE_NAME 128
#define RASSAPI_MAX_DEVICETYPE_NAME 16
#define RASSAPI_MAX_PARAM_KEY_SIZE 32
#define RASPRIV_NoCallback 0x01
#define RASPRIV_AdminSetCallback 0x02
#define RASPRIV_CallerSetCallback 0x04
#define RASPRIV_DialinPrivilege 0x08
#define RASPRIV_CallbackType 0x07
#define RAS_MODEM_OPERATIONAL 1
#define RAS_MODEM_NOT_RESPONDING 2
#define RAS_MODEM_HARDWARE_FAILURE 3
#define RAS_MODEM_INCORRECT_RESPONSE 4
#define RAS_MODEM_UNKNOWN 5
#define RAS_PORT_NON_OPERATIONAL 1
#define RAS_PORT_DISCONNECTED 2
#define RAS_PORT_CALLING_BACK 3
#define RAS_PORT_LISTENING 4
#define RAS_PORT_AUTHENTICATING 5
#define RAS_PORT_AUTHENTICATED 6
#define RAS_PORT_INITIALIZING 7
#define ParamNumber 0
#define ParamString 1
#define MEDIA_UNKNOWN 0
#define MEDIA_SERIAL 1
#define MEDIA_RAS10_SERIAL 2
#define MEDIA_X25 3
#define MEDIA_ISDN 4
#define USER_AUTHENTICATED 0x0001
#define MESSENGER_PRESENT 0x0002
#define PPP_CLIENT 0x0004
#define GATEWAY_ACTIVE 0x0008
#define REMOTE_LISTEN 0x0010
#define PORT_MULTILINKED 0x0020
#define RAS_IPADDRESSLEN 15
#define RAS_IPXADDRESSLEN 22
#define RAS_ATADDRESSLEN 32
#define RASDOWNLEVEL 10
#define RASADMIN_35 35
#define RASADMIN_CURRENT 40
#define RCD_SingleUser 0
#define RCD_AllUsers 0x00000001
#define RCD_Eap 0x00000002
#define RCD_Logon 0x00000004
#define CNLEN 15
#define LM20_CNLEN 15
#define DNLEN CNLEN
#define LM20_DNLEN LM20_CNLEN
#define UNCLEN (CNLEN+2)
#define LM20_UNCLEN (LM20_CNLEN+2)
#define NNLEN 80
#define LM20_NNLEN 12
#define RMLEN (UNCLEN+1+NNLEN)
#define LM20_RMLEN (LM20_UNCLEN+1+LM20_NNLEN)
#define SNLEN 80
#define LM20_SNLEN 15
#define STXTLEN 256
#define LM20_STXTLEN 63
#define PATHLEN 256
#define LM20_PATHLEN 256
#define DEVLEN 80
#define LM20_DEVLEN 8
#define EVLEN 16
#define UNLEN 256
#define LM20_UNLEN 20
#define GNLEN UNLEN
#define LM20_GNLEN LM20_UNLEN
#define PWLEN 256
#define LM20_PWLEN 14
#define SHPWLEN 8
#define CLTYPE_LEN 12
#define MAXCOMMENTSZ 256
#define LM20_MAXCOMMENTSZ 48
#define QNLEN NNLEN
#define LM20_QNLEN LM20_NNLEN
#define ALERTSZ 128
#define MAXDEVENTRIES 32
#define NETBIOS_NAME_LEN 16
#define MAX_PREFERRED_LENGTH ((DWORD) -1)
#define CRYPT_KEY_LEN 7
#define CRYPT_TXT_LEN 8
#define ENCRYPTED_PWLEN 16
#define SESSION_PWLEN 24
#define SESSION_CRYPT_KLEN 21
#define PARM_ERROR_UNKNOWN (-1)
#define PARM_ERROR_NONE 0
#define PARMNUM_BASE_INFOLEVEL 1000
#define MESSAGE_FILENAME "NETMSG"
#define OS2MSG_FILENAME "BASE"
#define HELP_MSG_FILENAME "NETH"
#define BACKUP_MSG_FILENAME "BAK.MSG"
#define PLATFORM_ID_DOS 300
#define PLATFORM_ID_OS2 400
#define PLATFORM_ID_NT 500
#define PLATFORM_ID_OSF 600
#define PLATFORM_ID_VMS 700
#define NERR_BASE 2100
#define MIN_LANMAN_MESSAGE_ID NERR_BASE
#define MAX_LANMAN_MESSAGE_ID 5799
#define NERR_Success 0
#define NERR_NetNotStarted (NERR_BASE+2)
#define NERR_UnknownServer (NERR_BASE+3)
#define NERR_ShareMem (NERR_BASE+4)
#define NERR_NoNetworkResource (NERR_BASE+5)
#define NERR_RemoteOnly (NERR_BASE+6)
#define NERR_DevNotRedirected (NERR_BASE+7)
#define NERR_ServerNotStarted (NERR_BASE+14)
#define NERR_ItemNotFound (NERR_BASE+15)
#define NERR_UnknownDevDir (NERR_BASE+16)
#define NERR_RedirectedPath (NERR_BASE+17)
#define NERR_DuplicateShare (NERR_BASE+18)
#define NERR_NoRoom (NERR_BASE+19)
#define NERR_TooManyItems (NERR_BASE+21)
#define NERR_InvalidMaxUsers (NERR_BASE+22)
#define NERR_BufTooSmall (NERR_BASE+23)
#define NERR_RemoteErr (NERR_BASE+27)
#define NERR_LanmanIniError (NERR_BASE+31)
#define NERR_NetworkError (NERR_BASE+36)
#define NERR_WkstaInconsistentState (NERR_BASE+37)
#define NERR_WkstaNotStarted (NERR_BASE+38)
#define NERR_BrowserNotStarted (NERR_BASE+39)
#define NERR_InternalError (NERR_BASE+40)
#define NERR_BadTransactConfig (NERR_BASE+41)
#define NERR_InvalidAPI (NERR_BASE+42)
#define NERR_BadEventName (NERR_BASE+43)
#define NERR_DupNameReboot (NERR_BASE+44)
#define NERR_CfgCompNotFound (NERR_BASE+46)
#define NERR_CfgParamNotFound (NERR_BASE+47)
#define NERR_LineTooLong (NERR_BASE+49)
#define NERR_QNotFound (NERR_BASE+50)
#define NERR_JobNotFound (NERR_BASE+51)
#define NERR_DestNotFound (NERR_BASE+52)
#define NERR_DestExists (NERR_BASE+53)
#define NERR_QExists (NERR_BASE+54)
#define NERR_QNoRoom (NERR_BASE+55)
#define NERR_JobNoRoom (NERR_BASE+56)
#define NERR_DestNoRoom (NERR_BASE+57)
#define NERR_DestIdle (NERR_BASE+58)
#define NERR_DestInvalidOp (NERR_BASE+59)
#define NERR_ProcNoRespond (NERR_BASE+60)
#define NERR_SpoolerNotLoaded (NERR_BASE+61)
#define NERR_DestInvalidState (NERR_BASE+62)
#define NERR_QInvalidState (NERR_BASE+63)
#define NERR_JobInvalidState (NERR_BASE+64)
#define NERR_SpoolNoMemory (NERR_BASE+65)
#define NERR_DriverNotFound (NERR_BASE+66)
#define NERR_DataTypeInvalid (NERR_BASE+67)
#define NERR_ProcNotFound (NERR_BASE+68)
#define NERR_ServiceTableLocked (NERR_BASE+80)
#define NERR_ServiceTableFull (NERR_BASE+81)
#define NERR_ServiceInstalled (NERR_BASE+82)
#define NERR_ServiceEntryLocked (NERR_BASE+83)
#define NERR_ServiceNotInstalled (NERR_BASE+84)
#define NERR_BadServiceName (NERR_BASE+85)
#define NERR_ServiceCtlTimeout (NERR_BASE+86)
#define NERR_ServiceCtlBusy (NERR_BASE+87)
#define NERR_BadServiceProgName (NERR_BASE+88)
#define NERR_ServiceNotCtrl (NERR_BASE+89)
#define NERR_ServiceKillProc (NERR_BASE+90)
#define NERR_ServiceCtlNotValid (NERR_BASE+91)
#define NERR_NotInDispatchTbl (NERR_BASE+92)
#define NERR_BadControlRecv (NERR_BASE+93)
#define NERR_ServiceNotStarting (NERR_BASE+94)
#define NERR_AlreadyLoggedOn (NERR_BASE+100)
#define NERR_NotLoggedOn (NERR_BASE+101)
#define NERR_BadUsername (NERR_BASE+102)
#define NERR_BadPassword (NERR_BASE+103)
#define NERR_UnableToAddName_W (NERR_BASE+104)
#define NERR_UnableToAddName_F (NERR_BASE+105)
#define NERR_UnableToDelName_W (NERR_BASE+106)
#define NERR_UnableToDelName_F (NERR_BASE+107)
#define NERR_LogonsPaused (NERR_BASE+109)
#define NERR_LogonServerConflict (NERR_BASE+110)
#define NERR_LogonNoUserPath (NERR_BASE+111)
#define NERR_LogonScriptError (NERR_BASE+112)
#define NERR_StandaloneLogon (NERR_BASE+114)
#define NERR_LogonServerNotFound (NERR_BASE+115)
#define NERR_LogonDomainExists (NERR_BASE+116)
#define NERR_NonValidatedLogon (NERR_BASE+117)
#define NERR_ACFNotFound (NERR_BASE+119)
#define NERR_GroupNotFound (NERR_BASE+120)
#define NERR_UserNotFound (NERR_BASE+121)
#define NERR_ResourceNotFound (NERR_BASE+122)
#define NERR_GroupExists (NERR_BASE+123)
#define NERR_UserExists (NERR_BASE+124)
#define NERR_ResourceExists (NERR_BASE+125)
#define NERR_NotPrimary (NERR_BASE+126)
#define NERR_ACFNotLoaded (NERR_BASE+127)
#define NERR_ACFNoRoom (NERR_BASE+128)
#define NERR_ACFFileIOFail (NERR_BASE+129)
#define NERR_ACFTooManyLists (NERR_BASE+130)
#define NERR_UserLogon (NERR_BASE+131)
#define NERR_ACFNoParent (NERR_BASE+132)
#define NERR_CanNotGrowSegment (NERR_BASE+133)
#define NERR_SpeGroupOp (NERR_BASE+134)
#define NERR_NotInCache (NERR_BASE+135)
#define NERR_UserInGroup (NERR_BASE+136)
#define NERR_UserNotInGroup (NERR_BASE+137)
#define NERR_AccountUndefined (NERR_BASE+138)
#define NERR_AccountExpired (NERR_BASE+139)
#define NERR_InvalidWorkstation (NERR_BASE+140)
#define NERR_InvalidLogonHours (NERR_BASE+141)
#define NERR_PasswordExpired (NERR_BASE+142)
#define NERR_PasswordCantChange (NERR_BASE+143)
#define NERR_PasswordHistConflict (NERR_BASE+144)
#define NERR_PasswordTooShort (NERR_BASE+145)
#define NERR_PasswordTooRecent (NERR_BASE+146)
#define NERR_InvalidDatabase (NERR_BASE+147)
#define NERR_DatabaseUpToDate (NERR_BASE+148)
#define NERR_SyncRequired (NERR_BASE+149)
#define NERR_UseNotFound (NERR_BASE+150)
#define NERR_BadAsgType (NERR_BASE+151)
#define NERR_DeviceIsShared (NERR_BASE+152)
#define NERR_NoComputerName (NERR_BASE+170)
#define NERR_MsgAlreadyStarted (NERR_BASE+171)
#define NERR_MsgInitFailed (NERR_BASE+172)
#define NERR_NameNotFound (NERR_BASE+173)
#define NERR_AlreadyForwarded (NERR_BASE+174)
#define NERR_AddForwarded (NERR_BASE+175)
#define NERR_AlreadyExists (NERR_BASE+176)
#define NERR_TooManyNames (NERR_BASE+177)
#define NERR_DelComputerName (NERR_BASE+178)
#define NERR_LocalForward (NERR_BASE+179)
#define NERR_GrpMsgProcessor (NERR_BASE+180)
#define NERR_PausedRemote (NERR_BASE+181)
#define NERR_BadReceive (NERR_BASE+182)
#define NERR_NameInUse (NERR_BASE+183)
#define NERR_MsgNotStarted (NERR_BASE+184)
#define NERR_NotLocalName (NERR_BASE+185)
#define NERR_NoForwardName (NERR_BASE+186)
#define NERR_RemoteFull (NERR_BASE+187)
#define NERR_NameNotForwarded (NERR_BASE+188)
#define NERR_TruncatedBroadcast (NERR_BASE+189)
#define NERR_InvalidDevice (NERR_BASE+194)
#define NERR_WriteFault (NERR_BASE+195)
#define NERR_DuplicateName (NERR_BASE+197)
#define NERR_DeleteLater (NERR_BASE+198)
#define NERR_IncompleteDel (NERR_BASE+199)
#define NERR_MultipleNets (NERR_BASE+200)
#define NERR_NetNameNotFound (NERR_BASE+210)
#define NERR_DeviceNotShared (NERR_BASE+211)
#define NERR_ClientNameNotFound (NERR_BASE+212)
#define NERR_FileIdNotFound (NERR_BASE+214)
#define NERR_ExecFailure (NERR_BASE+215)
#define NERR_TmpFile (NERR_BASE+216)
#define NERR_TooMuchData (NERR_BASE+217)
#define NERR_DeviceShareConflict (NERR_BASE+218)
#define NERR_BrowserTableIncomplete (NERR_BASE+219)
#define NERR_NotLocalDomain (NERR_BASE+220)
#define NERR_IsDfsShare (NERR_BASE+221)
#define NERR_DevInvalidOpCode (NERR_BASE+231)
#define NERR_DevNotFound (NERR_BASE+232)
#define NERR_DevNotOpen (NERR_BASE+233)
#define NERR_BadQueueDevString (NERR_BASE+234)
#define NERR_BadQueuePriority (NERR_BASE+235)
#define NERR_NoCommDevs (NERR_BASE+237)
#define NERR_QueueNotFound (NERR_BASE+238)
#define NERR_BadDevString (NERR_BASE+240)
#define NERR_BadDev (NERR_BASE+241)
#define NERR_InUseBySpooler (NERR_BASE+242)
#define NERR_CommDevInUse (NERR_BASE+243)
#define NERR_InvalidComputer (NERR_BASE+251)
#define NERR_MaxLenExceeded (NERR_BASE+254)
#define NERR_BadComponent (NERR_BASE+256)
#define NERR_CantType (NERR_BASE+257)
#define NERR_TooManyEntries (NERR_BASE+262)
#define NERR_ProfileFileTooBig (NERR_BASE+270)
#define NERR_ProfileOffset (NERR_BASE+271)
#define NERR_ProfileCleanup (NERR_BASE+272)
#define NERR_ProfileUnknownCmd (NERR_BASE+273)
#define NERR_ProfileLoadErr (NERR_BASE+274)
#define NERR_ProfileSaveErr (NERR_BASE+275)
#define NERR_LogOverflow (NERR_BASE+277)
#define NERR_LogFileChanged (NERR_BASE+278)
#define NERR_LogFileCorrupt (NERR_BASE+279)
#define NERR_SourceIsDir (NERR_BASE+280)
#define NERR_BadSource (NERR_BASE+281)
#define NERR_BadDest (NERR_BASE+282)
#define NERR_DifferentServers (NERR_BASE+283)
#define NERR_RunSrvPaused (NERR_BASE+285)
#define NERR_ErrCommRunSrv (NERR_BASE+289)
#define NERR_ErrorExecingGhost (NERR_BASE+291)
#define NERR_ShareNotFound (NERR_BASE+292)
#define NERR_InvalidLana (NERR_BASE+300)
#define NERR_OpenFiles (NERR_BASE+301)
#define NERR_ActiveConns (NERR_BASE+302)
#define NERR_BadPasswordCore (NERR_BASE+303)
#define NERR_DevInUse (NERR_BASE+304)
#define NERR_LocalDrive (NERR_BASE+305)
#define NERR_AlertExists (NERR_BASE+330)
#define NERR_TooManyAlerts (NERR_BASE+331)
#define NERR_NoSuchAlert (NERR_BASE+332)
#define NERR_BadRecipient (NERR_BASE+333)
#define NERR_AcctLimitExceeded (NERR_BASE+334)
#define NERR_InvalidLogSeek (NERR_BASE+340)
#define NERR_BadUasConfig (NERR_BASE+350)
#define NERR_InvalidUASOp (NERR_BASE+351)
#define NERR_LastAdmin (NERR_BASE+352)
#define NERR_DCNotFound (NERR_BASE+353)
#define NERR_LogonTrackingError (NERR_BASE+354)
#define NERR_NetlogonNotStarted (NERR_BASE+355)
#define NERR_CanNotGrowUASFile (NERR_BASE+356)
#define NERR_TimeDiffAtDC (NERR_BASE+357)
#define NERR_PasswordMismatch (NERR_BASE+358)
#define NERR_NoSuchServer (NERR_BASE+360)
#define NERR_NoSuchSession (NERR_BASE+361)
#define NERR_NoSuchConnection (NERR_BASE+362)
#define NERR_TooManyServers (NERR_BASE+363)
#define NERR_TooManySessions (NERR_BASE+364)
#define NERR_TooManyConnections (NERR_BASE+365)
#define NERR_TooManyFiles (NERR_BASE+366)
#define NERR_NoAlternateServers (NERR_BASE+367)
#define NERR_TryDownLevel (NERR_BASE+370)
#define NERR_UPSDriverNotStarted (NERR_BASE+380)
#define NERR_UPSInvalidConfig (NERR_BASE+381)
#define NERR_UPSInvalidCommPort (NERR_BASE+382)
#define NERR_UPSSignalAsserted (NERR_BASE+383)
#define NERR_UPSShutdownFailed (NERR_BASE+384)
#define NERR_BadDosRetCode (NERR_BASE+400)
#define NERR_ProgNeedsExtraMem (NERR_BASE+401)
#define NERR_BadDosFunction (NERR_BASE+402)
#define NERR_RemoteBootFailed (NERR_BASE+403)
#define NERR_BadFileCheckSum (NERR_BASE+404)
#define NERR_NoRplBootSystem (NERR_BASE+405)
#define NERR_RplLoadrNetBiosErr (NERR_BASE+406)
#define NERR_RplLoadrDiskErr (NERR_BASE+407)
#define NERR_ImageParamErr (NERR_BASE+408)
#define NERR_TooManyImageParams (NERR_BASE+409)
#define NERR_NonDosFloppyUsed (NERR_BASE+410)
#define NERR_RplBootRestart (NERR_BASE+411)
#define NERR_RplSrvrCallFailed (NERR_BASE+412)
#define NERR_CantConnectRplSrvr (NERR_BASE+413)
#define NERR_CantOpenImageFile (NERR_BASE+414)
#define NERR_CallingRplSrvr (NERR_BASE+415)
#define NERR_StartingRplBoot (NERR_BASE+416)
#define NERR_RplBootServiceTerm (NERR_BASE+417)
#define NERR_RplBootStartFailed (NERR_BASE+418)
#define NERR_RPL_CONNECTED (NERR_BASE+419)
#define NERR_BrowserConfiguredToNotRun (NERR_BASE+450)
#define NERR_RplNoAdaptersStarted (NERR_BASE+510)
#define NERR_RplBadRegistry (NERR_BASE+511)
#define NERR_RplBadDatabase (NERR_BASE+512)
#define NERR_RplRplfilesShare (NERR_BASE+513)
#define NERR_RplNotRplServer (NERR_BASE+514)
#define NERR_RplCannotEnum (NERR_BASE+515)
#define NERR_RplWkstaInfoCorrupted (NERR_BASE+516)
#define NERR_RplWkstaNotFound (NERR_BASE+517)
#define NERR_RplWkstaNameUnavailable (NERR_BASE+518)
#define NERR_RplProfileInfoCorrupted (NERR_BASE+519)
#define NERR_RplProfileNotFound (NERR_BASE+520)
#define NERR_RplProfileNameUnavailable (NERR_BASE+521)
#define NERR_RplProfileNotEmpty (NERR_BASE+522)
#define NERR_RplConfigInfoCorrupted (NERR_BASE+523)
#define NERR_RplConfigNotFound (NERR_BASE+524)
#define NERR_RplAdapterInfoCorrupted (NERR_BASE+525)
#define NERR_RplInternal (NERR_BASE+526)
#define NERR_RplVendorInfoCorrupted (NERR_BASE+527)
#define NERR_RplBootInfoCorrupted (NERR_BASE+528)
#define NERR_RplWkstaNeedsUserAcct (NERR_BASE+529)
#define NERR_RplNeedsRPLUSERAcct (NERR_BASE+530)
#define NERR_RplBootNotFound (NERR_BASE+531)
#define NERR_RplIncompatibleProfile (NERR_BASE+532)
#define NERR_RplAdapterNameUnavailable (NERR_BASE+533)
#define NERR_RplConfigNotEmpty (NERR_BASE+534)
#define NERR_RplBootInUse (NERR_BASE+535)
#define NERR_RplBackupDatabase (NERR_BASE+536)
#define NERR_RplAdapterNotFound (NERR_BASE+537)
#define NERR_RplVendorNotFound (NERR_BASE+538)
#define NERR_RplVendorNameUnavailable (NERR_BASE+539)
#define NERR_RplBootNameUnavailable (NERR_BASE+540)
#define NERR_RplConfigNameUnavailable (NERR_BASE+541)
#define NERR_DfsInternalCorruption (NERR_BASE+560)
#define NERR_DfsVolumeDataCorrupt (NERR_BASE+561)
#define NERR_DfsNoSuchVolume (NERR_BASE+562)
#define NERR_DfsVolumeAlreadyExists (NERR_BASE+563)
#define NERR_DfsAlreadyShared (NERR_BASE+564)
#define NERR_DfsNoSuchShare (NERR_BASE+565)
#define NERR_DfsNotALeafVolume (NERR_BASE+566)
#define NERR_DfsLeafVolume (NERR_BASE+567)
#define NERR_DfsVolumeHasMultipleServers (NERR_BASE+568)
#define NERR_DfsCantCreateJunctionPoint (NERR_BASE+569)
#define NERR_DfsServerNotDfsAware (NERR_BASE+570)
#define NERR_DfsBadRenamePath (NERR_BASE+571)
#define NERR_DfsVolumeIsOffline (NERR_BASE+572)
#define NERR_DfsInternalError (NERR_BASE+590)
#define MAX_NERR (NERR_BASE+899)
#define cchTextLimitDefault 32767
#define WM_CONTEXTME 0x007B
#define EM_CANPASTE (WM_USER + 50)
#define EM_DISPLAYBAND (WM_USER + 51)
#define EM_EXGETSEL (WM_USER + 52)
#define EM_EXLIMITTEXT (WM_USER + 53)
#define EM_EXLINEFROMCHAR (WM_USER + 54)
#define EM_EXSETSEL (WM_USER + 55)
#define EM_FINDTEXT (WM_USER + 56)
#define EM_FORMATRANGE (WM_USER + 57)
#define EM_GETCHARFORMAT (WM_USER + 58)
#define EM_GETEVENTMASK (WM_USER + 59)
#define EM_GETOLEINTERFACE (WM_USER + 60)
#define EM_GETPARAFORMAT (WM_USER + 61)
#define EM_GETSELTEXT (WM_USER + 62)
#define EM_HIDESELECTION (WM_USER + 63)
#define EM_PASTESPECIAL (WM_USER + 64)
#define EM_REQUESTRESIZE (WM_USER + 65)
#define EM_SELECTIONTYPE (WM_USER + 66)
#define EM_SETBKGNDCOLOR (WM_USER + 67)
#define EM_SETCHARFORMAT (WM_USER + 68)
#define EM_SETEVENTMASK (WM_USER + 69)
#define EM_SETOLECALLBACK (WM_USER + 70)
#define EM_SETPARAFORMAT (WM_USER + 71)
#define EM_SETTARGETDEVICE (WM_USER + 72)
#define EM_STREAMIN (WM_USER + 73)
#define EM_STREAMOUT (WM_USER + 74)
#define EM_GETTEXTRANGE (WM_USER + 75)
#define EM_FINDWORDBREAK (WM_USER + 76)
#define EM_SETOPTIONS (WM_USER + 77)
#define EM_GETOPTIONS (WM_USER + 78)
#define EM_FINDTEXTEX (WM_USER + 79)
#define EM_GETWORDBREAKPROCEX (WM_USER + 80)
#define EM_SETWORDBREAKPROCEX (WM_USER + 81)
#define EM_SHOWSCROLLBAR (WM_USER + 96)
#define EM_SETTEXTEX (WM_USER + 97)
#define EM_SETPUNCTUATION (WM_USER + 100)
#define EM_GETPUNCTUATION (WM_USER + 101)
#define EM_SETWORDWRAPMODE (WM_USER + 102)
#define EM_GETWORDWRAPMODE (WM_USER + 103)
#define EM_SETIMECOLOR (WM_USER + 104)
#define EM_GETIMECOLOR (WM_USER + 105)
#define EM_SETIMEOPTIONS (WM_USER + 106)
#define EM_GETIMEOPTIONS (WM_USER + 107)
#define EM_CONVPOSITION (WM_USER + 108)
#define EM_SETLANGOPTIONS (WM_USER + 120)
#define EM_GETLANGOPTIONS (WM_USER + 121)
#define EM_GETIMECOMPMODE (WM_USER + 122)
#define EM_FINDTEXTW (WM_USER + 123)
#define EM_FINDTEXTEXW ( WM_USER + 124)
#define EM_RECONVERSION (WM_USER + 125)
#define EM_SETIMEMODEBIAS (WM_USER + 126)
#define EM_GETIMEMODEBIAS (WM_USER + 127)
#define EM_SETBIDIOPTIONS (WM_USER + 200)
#define EM_GETBIDIOPTIONS (WM_USER + 201)
#define EM_SETTYPOGRAPHYOPTIONS (WM_USER + 202)
#define EM_GETTYPOGRAPHYOPTIONS (WM_USER + 203)
#define EM_SETEDITSTYLE (WM_USER + 204)
#define EM_GETEDITSTYLE (WM_USER + 205)
#define SES_EMULATESYSEDIT 1
#define SES_BEEPONMAXTEXT 2
#define SES_EXTENDBACKCOLOR 4
#define SES_MAPCPS 8
#define SES_EMULATE10 16
#define SES_USECRLF 32
#define SES_USEAIMM 64
#define SES_NOIME 128
#define SES_ALLOWBEEPS 256
#define SES_UPPERCASE 512
#define SES_LOWERCASE 1024
#define SES_NOINPUTSEQUENCECHK 2048
#define SES_BIDI 4096
#define SES_SCROLLONKILLFOCUS 8192
#define SES_XLTCRCRLFTOCR 16384
#define SES_DRAFTMODE 32768
#define SES_USECTF 0x0010000
#define SES_HIDEGRIDLINES 0x0020000
#define SES_USEATFONT 0x0040000
#define SES_CUSTOMLOOK 0x0080000
#define SES_LBSCROLLNOTIFY 0x0100000
#define SES_CTFALLOWEMBED 0x0200000
#define SES_CTFALLOWSMARTTAG 0x0400000
#define SES_CTFALLOWPROOFING 0x0800000
#define IMF_AUTOKEYBOARD 0x0001
#define IMF_AUTOFONT 0x0002
#define IMF_IMECANCELCOMPLETE 0x0004
#define IMF_IMEALWAYSSENDNOTIFY 0x0008
#define IMF_AUTOFONTSIZEADJUST 0x0010
#define IMF_UIFONTS 0x0020
#define IMF_DUALFONT 0x0080
#define ICM_NOTOPEN 0x0000
#define ICM_LEVEL3 0x0001
#define ICM_LEVEL2 0x0002
#define ICM_LEVEL2_5 0x0003
#define ICM_LEVEL2_SUI 0x0004
#define ICM_CTF 0x0005
#define TO_ADVANCEDTYPOGRAPHY 1
#define TO_SIMPLELINEBREAK 2
#define TO_DISABLECUSTOMTEXTOUT 4
#define TO_ADVANCEDLAYOUT 8
#define EM_OUTLINE (WM_USER + 220)
#define EM_GETSCROLLPOS (WM_USER + 221)
#define EM_SETSCROLLPOS (WM_USER + 222)
#define EM_SETFONTSIZE (WM_USER + 223)
#define EM_GETZOOM (WM_USER + 224)
#define EM_SETZOOM (WM_USER + 225)
#define EM_GETVIEWKIND (WM_USER + 226)
#define EM_SETVIEWKIND (WM_USER + 227)
#define EM_GETPAGE (WM_USER + 228)
#define EM_SETPAGE (WM_USER + 229)
#define EM_GETHYPHENATEINFO (WM_USER + 230)
#define EM_SETHYPHENATEINFO (WM_USER + 231)
#define EM_GETPAGEROTATE (WM_USER + 235)
#define EM_SETPAGEROTATE (WM_USER + 236)
#define EM_GETCTFMODEBIAS (WM_USER + 237)
#define EM_SETCTFMODEBIAS (WM_USER + 238)
#define EM_GETCTFOPENSTATUS (WM_USER + 240)
#define EM_SETCTFOPENSTATUS (WM_USER + 241)
#define EM_GETIMECOMPTEXT (WM_USER + 242)
#define EM_ISIME (WM_USER + 243)
#define EM_GETIMEPROPERTY (WM_USER + 244)
#define EM_GETQUERYRTFOBJ (WM_USER + 269)
#define EM_SETQUERYRTFOBJ (WM_USER + 270)
#define EPR_0 0
#define EPR_270 1
#define EPR_180 2
#define EPR_90 3
#define CTFMODEBIAS_DEFAULT 0x0000
#define CTFMODEBIAS_FILENAME 0x0001
#define CTFMODEBIAS_NAME 0x0002
#define CTFMODEBIAS_READING 0x0003
#define CTFMODEBIAS_DATETIME 0x0004
#define CTFMODEBIAS_CONVERSATION 0x0005
#define CTFMODEBIAS_NUMERIC 0x0006
#define CTFMODEBIAS_HIRAGANA 0x0007
#define CTFMODEBIAS_KATAKANA 0x0008
#define CTFMODEBIAS_HANGUL 0x0009
#define CTFMODEBIAS_HALFWIDTHKATAKANA 0x000A
#define CTFMODEBIAS_FULLWIDTHALPHANUMERIC 0x000B
#define CTFMODEBIAS_HALFWIDTHALPHANUMERIC 0x000C
#define IMF_SMODE_PLAURALCLAUSE 0x0001
#define IMF_SMODE_NONE 0x0002
#define EMO_EXIT 0
#define EMO_ENTER 1
#define EMO_PROMOTE 2
#define EMO_EXPAND 3
#define EMO_MOVESELECTION 4
#define EMO_GETVIEWMODE 5
#define EMO_EXPANDSELECTION 0
#define EMO_EXPANDDOCUMENT 1
#define VM_NORMAL 4
#define VM_OUTLINE 2
#define VM_PAGE 9
#define EN_MSGFILTER 0x0700
#define EN_REQUESTRESIZE 0x0701
#define EN_SELCHANGE 0x0702
#define EN_DROPFILES 0x0703
#define EN_PROTECTED 0x0704
#define EN_CORRECTTEXT 0x0705
#define EN_STOPNOUNDO 0x0706
#define EN_IMECHANGE 0x0707
#define EN_SAVECLIPBOARD 0x0708
#define EN_OLEOPFAILED 0x0709
#define EN_OBJECTPOSITIONS 0x070a
#define EN_LINK 0x070b
#define EN_DRAGDROPDONE 0x070c
#define EN_PARAGRAPHEXPANDED 0x070d
#define EN_PAGECHANGE 0x070e
#define EN_LOWFIRTF 0x070f
#define EN_ALIGNLTR 0x0710
#define EN_ALIGNRTL 0x0711
#define ENM_NONE 0x00000000
#define ENM_CHANGE 0x00000001
#define ENM_UPDATE 0x00000002
#define ENM_SCROLL 0x00000004
#define ENM_SCROLLEVENTS 0x00000008
#define ENM_DRAGDROPDONE 0x00000010
#define ENM_PARAGRAPHEXPANDED 0x00000020
#define ENM_PAGECHANGE 0x00000040
#define ENM_KEYEVENTS 0x00010000
#define ENM_MOUSEEVENTS 0x00020000
#define ENM_REQUESTRESIZE 0x00040000
#define ENM_SELCHANGE 0x00080000
#define ENM_DROPFILES 0x00100000
#define ENM_PROTECTED 0x00200000
#define ENM_CORRECTTEXT 0x00400000
#define ENM_IMECHANGE 0x00800000
#define ENM_LANGCHANGE 0x01000000
#define ENM_OBJECTPOSITIONS 0x02000000
#define ENM_LINK 0x04000000
#define ENM_LOWFIRTF 0x08000000
#define ES_SAVESEL 0x00008000
#define ES_SUNKEN 0x00004000
#define ES_DISABLENOSCROLL 0x00002000
#define ES_SELECTIONBAR 0x01000000
#define ES_NOOLEDRAGDROP 0x00000008
#define ES_EX_NOCALLOLEINIT 0x01000000
#define ES_VERTICAL 0x00400000
#define ES_NOIME 0x00080000
#define ES_SELFIME 0x00040000
#define ECO_AUTOWORDSELECTION 0x00000001
#define ECO_AUTOVSCROLL 0x00000040
#define ECO_AUTOHSCROLL 0x00000080
#define ECO_NOHIDESEL 0x00000100
#define ECO_READONLY 0x00000800
#define ECO_WANTRETURN 0x00001000
#define ECO_SAVESEL 0x00008000
#define ECO_SELECTIONBAR 0x01000000
#define ECO_VERTICAL 0x00400000
#define ECOOP_SET 0x0001
#define ECOOP_OR 0x0002
#define ECOOP_AND 0x0003
#define ECOOP_XOR 0x0004
#define WB_CLASSIFY 3
#define WB_MOVEWORDLEFT 4
#define WB_MOVEWORDRIGHT 5
#define WB_LEFTBREAK 6
#define WB_RIGHTBREAK 7
#define WB_MOVEWORDPREV 4
#define WB_MOVEWORDNEXT 5
#define WB_PREVBREAK 6
#define WB_NEXTBREAK 7
#define PC_FOLLOWING 1
#define PC_LEADING 2
#define PC_OVERFLOW 3
#define PC_DELIMITER 4
#define WBF_WORDWRAP 0x010
#define WBF_WORDBREAK 0x020
#define WBF_OVERFLOW 0x040
#define WBF_LEVEL1 0x080
#define WBF_LEVEL2 0x100
#define WBF_CUSTOM 0x200
#define IMF_FORCENONE 0x0001
#define IMF_FORCEENABLE 0x0002
#define IMF_FORCEDISABLE 0x0004
#define IMF_CLOSESTATUSWINDOW 0x0008
#define IMF_VERTICAL 0x0020
#define IMF_FORCEACTIVE 0x0040
#define IMF_FORCEINACTIVE 0x0080
#define IMF_FORCEREMEMBER 0x0100
#define IMF_MULTIPLEEDIT 0x0400
#define WBF_CLASS BYTE(_CAST,0x0F)
#define WBF_ISWHITE BYTE(_CAST,0x10)
#define WBF_BREAKLINE BYTE(_CAST,0x20)
#define WBF_BREAKAFTER BYTE(_CAST,0x40)
#define CFM_BOLD 0x00000001
#define CFM_ITALIC 0x00000002
#define CFM_UNDERLINE 0x00000004
#define CFM_STRIKEOUT 0x00000008
#define CFM_PROTECTED 0x00000010
#define CFM_LINK 0x00000020
#define CFM_SIZE 0x80000000L
#define CFM_COLOR 0x40000000L
#define CFM_FACE 0x20000000L
#define CFM_OFFSET 0x10000000L
#define CFM_CHARSET 0x08000000L
#define CFE_BOLD 0x0001
#define CFE_ITALIC 0x0002
#define CFE_UNDERLINE 0x0004
#define CFE_STRIKEOUT 0x0008
#define CFE_PROTECTED 0x0010
#define CFE_LINK 0x0020
#define CFE_AUTOCOLOR 0x40000000
#define CFM_SMALLCAPS 0x0040
#define CFM_ALLCAPS 0x0080
#define CFM_HIDDEN 0x0100
#define CFM_OUTLINE 0x0200
#define CFM_SHADOW 0x0400
#define CFM_EMBOSS 0x0800
#define CFM_IMPRINT 0x1000
#define CFM_DISABLED 0x2000
#define CFM_REVISED 0x4000
#define CFM_BACKCOLOR 0x04000000L
#define CFM_LCID 0x02000000L
#define CFM_UNDERLINETYPE 0x00800000L 
#define CFM_WEIGHT 0x00400000L
#define CFM_SPACING 0x00200000L 
#define CFM_KERNING 0x00100000L 
#define CFM_STYLE 0x00080000L 
#define CFM_ANIMATION 0x00040000L 
#define CFM_REVAUTHOR 0x00008000L
#define CFE_SUBSCRIPT 0x00010000
#define CFE_SUPERSCRIPT 0x00020000
#define CFM_SUBSCRIPT CFE_SUBSCRIPT | CFE_SUPERSCRIPT
#define CFM_SUPERSCRIPT CFM_SUBSCRIPT
#define CFM_EFFECTS (CFM_BOLD | CFM_ITALIC | CFM_UNDERLINE | CFM_COLOR | CFM_STRIKEOUT | CFE_PROTECTED | CFM_LINK)
#define CFM_ALL (CFM_EFFECTS | CFM_SIZE | CFM_FACE | CFM_OFFSET | CFM_CHARSET)
#define CFM_EFFECTS2 (CFM_EFFECTS | CFM_DISABLED | CFM_SMALLCAPS | CFM_ALLCAPS | CFM_HIDDEN | CFM_OUTLINE | CFM_SHADOW | CFM_EMBOSS | CFM_IMPRINT | CFM_DISABLED | CFM_REVISED | CFM_SUBSCRIPT | CFM_SUPERSCRIPT | CFM_BACKCOLOR)
#define CFM_ALL2 (CFM_ALL | CFM_EFFECTS2 | CFM_BACKCOLOR | CFM_LCID | CFM_UNDERLINETYPE | CFM_WEIGHT | CFM_REVAUTHOR | CFM_SPACING | CFM_KERNING | CFM_STYLE | CFM_ANIMATION)
#define CFE_SMALLCAPS CFM_SMALLCAPS
#define CFE_ALLCAPS CFM_ALLCAPS
#define CFE_HIDDEN CFM_HIDDEN
#define CFE_OUTLINE CFM_OUTLINE
#define CFE_SHADOW CFM_SHADOW
#define CFE_EMBOSS CFM_EMBOSS
#define CFE_IMPRINT CFM_IMPRINT
#define CFE_DISABLED CFM_DISABLED
#define CFE_REVISED CFM_REVISED
#define CFE_AUTOBACKCOLOR CFM_BACKCOLOR
#define CFU_CF1UNDERLINE 0xFF
#define CFU_INVERT 0xFE
#define CFU_UNDERLINETHICKLONGDASH 18
#define CFU_UNDERLINETHICKDOTTED 17
#define CFU_UNDERLINETHICKDASHDOTDOT 16
#define CFU_UNDERLINETHICKDASHDOT 15
#define CFU_UNDERLINETHICKDASH 14
#define CFU_UNDERLINELONGDASH 13
#define CFU_UNDERLINEHEAVYWAVE 12
#define CFU_UNDERLINEDOUBLEWAVE 11
#define CFU_UNDERLINEHAIRLINE 10
#define CFU_UNDERLINETHICK 9
#define CFU_UNDERLINEWAVE 8
#define CFU_UNDERLINEDASHDOTDOT 7
#define CFU_UNDERLINEDASHDOT 6
#define CFU_UNDERLINEDASH 5
#define CFU_UNDERLINEDOTTED 4
#define CFU_UNDERLINEDOUBLE 3
#define CFU_UNDERLINEWORD 2
#define CFU_UNDERLINE 1
#define CFU_UNDERLINENONE 0
#define yHeightCharPtsMost 1638
#define SCF_SELECTION 0x0001
#define SCF_WORD 0x0002
#define SCF_DEFAULT 0x0000
#define SCF_ALL 0x0004
#define SCF_USEUIRULES 0x0008
#define SCF_ASSOCIATEFONT 0x0010
#define SCF_NOKBUPDATE 0x0020
#define SCF_ASSOCIATEFONT2 0x0040
#define SF_TEXT 0x0001
#define SF_RTF 0x0002
#define SF_RTFNOOBJS 0x0003
#define SF_TEXTIZED 0x0004
#define SF_UNICODE 0x0010
#define SF_USECODEPAGE 0x0020
#define SF_NCRFORNONASCII 0x40
#define SFF_WRITEXTRAPAR 0x80
#define SFF_SELECTION 0x8000
#define SFF_PLAINRTF 0x4000
#define SFF_PERSISTVIEWSCALE 0x2000
#define SFF_KEEPDOCINFO 0x1000
#define SFF_PWD 0x0800
#define SF_RTFVAL 0x0700
#define MAX_TAB_STOPS 32
#define lDefaultTab 720
#define PFM_STARTINDENT 0x00000001
#define PFM_RIGHTINDENT 0x00000002
#define PFM_OFFSET 0x00000004
#define PFM_ALIGNMENT 0x00000008
#define PFM_TABSTOPS 0x00000010
#define PFM_NUMBERING 0x00000020
#define PFM_OFFSETINDENT 0x80000000
#define PFM_SPACEBEFORE 0x00000040L
#define PFM_SPACEAFTER 0x00000080L
#define PFM_LINESPACING 0x00000100L
#define PFM_STYLE 0x00000400L
#define PFM_BORDER 0x00000800L 
#define PFM_SHADING 0x00001000L 
#define PFM_NUMBERINGSTYLE 0x00002000L 
#define PFM_NUMBERINGTAB 0x00004000L 
#define PFM_NUMBERINGSTART 0x00008000L 
#define PFM_DIR 0x00010000L
#define PFM_RTLPARA 0x00010000L 
#define PFM_KEEP 0x00020000L 
#define PFM_KEEPNEXT 0x00040000L 
#define PFM_PAGEBREAKBEFORE 0x00080000L 
#define PFM_NOLINENUMBER 0x00100000L 
#define PFM_NOWIDOWCONTROL 0x00200000L 
#define PFM_DONOTHYPHEN 0x00400000L 
#define PFM_SIDEBYSIDE 0x00800000L 
#define PFM_TABLE 0xc0000000L 
#define PFM_TABLE_RE3 0x40000000
#define PFM_TEXTWRAPPINGBREAK 0x20000000
#define PFM_TABLEROWDELIMITER 0x10000000
#define PFM_COLLAPSED 0x01000000
#define PFM_OUTLINELEVEL 0x02000000
#define PFM_BOX 0x04000000
#define PFM_RESERVED2 0x08000000
#define PFM_ALL (PFM_STARTINDENT | PFM_RIGHTINDENT | PFM_OFFSET | PFM_ALIGNMENT | PFM_TABSTOPS | PFM_NUMBERING | PFM_OFFSETINDENT| PFM_RTLPARA)
#define PFM_EFFECTS (PFM_RTLPARA | PFM_KEEP | PFM_KEEPNEXT | PFM_TABLE | PFM_PAGEBREAKBEFORE | PFM_NOLINENUMBER | PFM_NOWIDOWCONTROL | PFM_DONOTHYPHEN | PFM_SIDEBYSIDE | PFM_TABLE | PFM_TABLEROWDELIMITER)
#define PFM_ALL2 (PFM_ALL | PFM_EFFECTS | PFM_SPACEBEFORE | PFM_SPACEAFTER | PFM_LINESPACING | PFM_STYLE | PFM_SHADING | PFM_BORDER | PFM_NUMBERINGTAB | PFM_NUMBERINGSTART | PFM_NUMBERINGSTYLE)
#define PFE_RTLPARA (PFM_RTLPARA >> 16)
#define PFE_KEEP (PFM_KEEP >> 16)
#define PFE_KEEPNEXT (PFM_KEEPNEXT >> 16)
#define PFE_PAGEBREAKBEFORE (PFM_PAGEBREAKBEFORE >> 16)
#define PFE_NOLINENUMBER (PFM_NOLINENUMBER >> 16)
#define PFE_NOWIDOWCONTROL (PFM_NOWIDOWCONTROL >> 16)
#define PFE_SIDEBYSIDE (PFM_SIDEBYSIDE >> 16)
#define PFE_TEXTWRAPPINGBREAK (PFM_TEXTWRAPPINGBREAK>>16)
#define PFE_COLLAPSED (PFM_COLLAPSED >> 16)
#define PFE_BOX (PFM_BOX >> 16)
#define PFN_BULLET 1
#define PFN_ARABIC 2
#define PFN_LCLETTER 3
#define PFN_UCLETTER 4
#define PFN_LCROMAN 5
#define PFN_UCROMAN 6
#define PFNS_PAREN 0x000
#define PFNS_PARENS 0x100
#define PFNS_PERIOD 0x200
#define PFNS_PLAIN 0x300
#define PFNS_NONUMBER 0x400
#define PFNS_NEWNUMBER 0x8000
#define PFA_LEFT 0x0001
#define PFA_RIGHT 0x0002
#define PFA_CENTER 0x0003
#define PFA_JUSTIFY 4
#define PFA_FULL_INTERWORD 4
#define PFA_FULL_INTERLETTER 5
#define PFA_FULL_SCALED 6
#define PFA_FULL_GLYPHS 7
#define PFA_SNAP_GRID 8
#define SEL_EMPTY 0x0000
#define SEL_TEXT 0x0001
#define SEL_OBJECT 0x0002
#define SEL_MULTICHAR 0x0004
#define SEL_MULTIOBJECT 0x0008
#define GCM_RIGHTMOUSEDROP 0x8000
#define OLEOP_DOVERB 1
#define CF_RTF "Rich Text Format"
#define CF_RTFNOOBJS "Rich Text Format Without Objects"
#define CF_RETEXTOBJ "RichEdit Text and Objects"
#define PFE_TABLEROW 0xc000 
#define PFE_TABLECELLEND 0x8000 
#define PFE_TABLECELL 0x4000 
#define ABM_NEW 0x00000000
#define ABM_REMOVE 0x00000001
#define ABM_QUERYPOS 0x00000002
#define ABM_SETPOS 0x00000003
#define ABM_GETSTATE 0x00000004
#define ABM_GETTASKBARPOS 0x00000005
#define ABM_ACTIVATE 0x00000006
#define ABM_GETAUTOHIDEBAR 0x00000007
#define ABM_SETAUTOHIDEBAR 0x00000008
#define ABM_WINDOWPOSCHANGED 0x0000009
#define ABM_SETSTATE 0x0000000a
#define ABN_STATECHANGE 0x0000000
#define ABN_POSCHANGED 0x0000001
#define ABN_FULLSCREENAPP 0x0000002
#define ABN_WINDOWARRANGE 0x0000003
#define ABS_AUTOHIDE 0x0000001
#define ABS_ALWAYSONTOP 0x0000002
#define ABE_LEFT 0
#define ABE_TOP 1
#define ABE_RIGHT 2
#define ABE_BOTTOM 3
#define FO_MOVE 0x0001
#define FO_COPY 0x0002
#define FO_DELETE 0x0003
#define FO_RENAME 0x0004
#define FOF_MULTIDESTFILES 0x0001
#define FOF_CONFIRMMOUSE 0x0002
#define FOF_SILENT 0x0004
#define FOF_RENAMEONCOLLISION 0x0008
#define FOF_NOCONFIRMATION 0x0010
#define FOF_WANTMAPPINGHANDLE 0x0020
#define FOF_ALLOWUNDO 0x0040
#define FOF_FILESONLY 0x0080
#define FOF_SIMPLEPROGRESS 0x0100
#define FOF_NOCONFIRMMKDIR 0x0200
#define FOF_NOERRORUI 0x0400
#define FOF_NOCOPYSECURITYATTRIBS 0x0800
#define FOF_NORECURSION 0x1000
#define FOF_NO_CONNECTED_ELEMENTS 0x2000
#define FOF_WANTNUKEWARNING 0x4000
#define FOF_NORECURSEREPARSE 0x8000
#define PO_DELETE 0x0013
#define PO_RENAME 0x0014
#define PO_PORTCHANGE 0x0020
#define PO_REN_PORT 0x0034
#define SE_ERR_FNF 2
#define SE_ERR_PNF 3
#define SE_ERR_ACCESSDENIED 5
#define SE_ERR_OOM 8
#define SE_ERR_DLLNOTFOUND 32
#define SE_ERR_SHARE 26
#define SE_ERR_ASSOCINCOMPLETE 27
#define SE_ERR_DDETIMEOUT 28
#define SE_ERR_DDEFAIL 29
#define SE_ERR_DDEBUSY 30
#define SE_ERR_NOASSOC 31
#define SEE_MASK_CLASSNAME 0x00000001
#define SEE_MASK_CLASSKEY 0x00000003
#define SEE_MASK_IDLIST 0x00000004
#define SEE_MASK_INVOKEIDLIST 0x0000000c
#define SEE_MASK_ICON 0x00000010
#define SEE_MASK_HOTKEY 0x00000020
#define SEE_MASK_NOCLOSEPROCESS 0x00000040
#define SEE_MASK_CONNECTNETDRV 0x00000080
#define SEE_MASK_FLAG_DDEWAIT 0x00000100
#define SEE_MASK_DOENVSUBST 0x00000200
#define SEE_MASK_FLAG_NO_UI 0x00000400
#define SEE_MASK_UNICODE 0x00010000
#define SEE_MASK_NO_CONSOLE 0x00008000
#define SEE_MASK_ASYNCOK 0x00100000
#define SEE_MASK_HMONITOR 0x00200000
#define SEE_MASK_NOZONECHECKS 0x00800000
#define SEE_MASK_NOQUERYCLASSSTORE 0x01000000
#define SEE_MASK_WAITFORINPUTIDLE 0x02000000
#define SEE_MASK_FLAG_LOG_USAGE 0x04000000
#define NIN_BALLOONSHOW (WM_USER + 2)
#define NIN_BALLOONHIDE (WM_USER + 3)
#define NIN_BALLOONTIMEOUT (WM_USER + 4)
#define NIN_BALLOONUSERCLICK (WM_USER + 5)
#define NIM_ADD 0x00000000
#define NIM_MODIFY 0x00000001
#define NIM_DELETE 0x00000002
#define NIM_SETFOCUS 0x00000003
#define NIM_SETVERSION 0x00000004
#define NOTIFYICON_VERSION 0x00000003
#define NIF_MESSAGE 0x00000001
#define NIF_ICON 0x00000002
#define NIF_TIP 0x00000004
#define NIF_STATE 0x00000008
#define NIF_INFO 0x00000010
#define NIF_GUID 0x00000020
#define NIS_HIDDEN 0x00000001
#define NIS_SHAREDICON 0x00000002
#define NIIF_NONE 0x00
#define NIIF_INFO 0x01
#define NIIF_WARNING 0x02
#define NIIF_ERROR 0x03
#define NIIF_USER 0x00000004
#define NIIF_ICON_MASK 0x0000000F
#define NIIF_NOSOUND 0x00000010
#define SHGFI_ICON 0x00000100
#define SHGFI_DISPLAYNAME 0x00000200
#define SHGFI_TYPENAME 0x00000400
#define SHGFI_ATTRIBUTES 0x00000800
#define SHGFI_ICONLOCATION 0x00001000
#define SHGFI_EXETYPE 0x00002000
#define SHGFI_SYSICONINDEX 0x00004000
#define SHGFI_LINKOVERLAY 0x00008000
#define SHGFI_SELECTED 0x00010000
#define SHGFI_ATTR_SPECIFIED 0x00020000
#define SHGFI_LARGEICON 0x00000000
#define SHGFI_SMALLICON 0x00000001
#define SHGFI_OPENICON 0x00000002
#define SHGFI_SHELLICONSIZE 0x00000004
#define SHGFI_PIDL 0x00000008
#define SHGFI_USEFILEATTRIBUTES 0x00000010
#define SHGFI_ADDOVERLAYS 0x00000020
#define SHGFI_OVERLAYINDEX 0x00000040
#define SHGNLI_PIDL 0x00000001
#define SHGNLI_PREFIXNAME 0x00000002
#define SHGNLI_NOUNIQUE 0x00000004
#define SHGNLI_NOLNK 0x00000008
#define SHACF_DEFAULT 0x00000000
#define SHACF_FILESYSTEM 0x00000001
#define SHACF_URLALL 0x00000006
#define SHACF_URLHISTORY 0x00000002
#define SHACF_URLMRU 0x00000004
#define SHACF_USETAB 0x00000008
#define SHACF_FILESYS_ONLY 0x00000010
#define SHACF_FILESYS_DIRS 0x00000020
#define SHACF_AUTOSUGGEST_FORCE_ON 0x10000000
#define SHACF_AUTOSUGGEST_FORCE_OFF 0x20000000
#define SHACF_AUTOAPPEND_FORCE_ON 0x40000000
#define SHACF_AUTOAPPEND_FORCE_OFF 0x80000000
#define SHGFP_TYPE_CURRENT 0
#define SHGFP_TYPE_DEFAULT 1
#define CSIDL_DESKTOP 0x0000
#define CSIDL_INTERNET 0x0001
#define CSIDL_PROGRAMS 0x0002
#define CSIDL_CONTROLS 0x0003
#define CSIDL_PRINTERS 0x0004
#define CSIDL_PERSONAL 0x0005
#define CSIDL_FAVORITES 0x0006
#define CSIDL_STARTUP 0x0007
#define CSIDL_RECENT 0x0008
#define CSIDL_SENDTO 0x0009
#define CSIDL_BITBUCKET 0x000A
#define CSIDL_STARTMENU 0x000B
#define CSIDL_MYDOCUMENTS 0x000c
#define CSIDL_MYMUSIC 0x000d
#define CSIDL_MYVIDEO 0x000e
#define CSIDL_DESKTOPDIRECTORY 0x0010
#define CSIDL_DRIVES 0x0011
#define CSIDL_NETWORK 0x0012
#define CSIDL_NETHOOD 0x0013
#define CSIDL_FONTS 0x0014
#define CSIDL_TEMPLATES 0x0015
#define CSIDL_COMMON_STARTMENU 0x0016
#define CSIDL_COMMON_PROGRAMS 0x0017
#define CSIDL_COMMON_STARTUP 0x0018
#define CSIDL_COMMON_DESKTOPDIRECTORY 0x0019
#define CSIDL_APPDATA 0x001A
#define CSIDL_PRINTHOOD 0x001B
#define CSIDL_LOCAL_APPDATA 0x001C
#define CSIDL_ALTSTARTUP 0x001D
#define CSIDL_COMMON_ALTSTARTUP 0x001E
#define CSIDL_COMMON_FAVORITES 0x001F
#define CSIDL_INTERNET_CACHE 0x0020
#define CSIDL_COOKIES 0x0021
#define CSIDL_HISTORY 0x0022
#define CSIDL_COMMON_APPDATA 0x0023
#define CSIDL_WINDOWS 0x0024
#define CSIDL_SYSTEM 0x0025
#define CSIDL_PROGRAM_FILES 0x0026
#define CSIDL_MYPICTURES 0x0027
#define CSIDL_PROFILE 0x0028
#define CSIDL_SYSTEMX86 0x0029
#define CSIDL_PROGRAM_FILESX86 0x002a
#define CSIDL_PROGRAM_FILES_COMMON 0x002b
#define CSIDL_PROGRAM_FILES_COMMONX86 0x002c
#define CSIDL_COMMON_TEMPLATES 0x002d
#define CSIDL_COMMON_DOCUMENTS 0x002e
#define CSIDL_COMMON_ADMINTOOLS 0x002f
#define CSIDL_ADMINTOOLS 0x0030
#define CSIDL_CONNECTIONS 0x0031
#define CSIDL_COMMON_MUSIC 0x0035
#define CSIDL_COMMON_PICTURES 0x0036
#define CSIDL_COMMON_VIDEO 0x0037
#define CSIDL_RESOURCES 0x0038
#define CSIDL_RESOURCES_LOCALIZED 0x0039
#define CSIDL_COMMON_OEM_LINKS 0x003a
#define CSIDL_CDBURN_AREA 0x003b
#define CSIDL_COMPUTERSNEARME 0x003d
#define CSIDL_FLAG_CREATE 0x8000
#define CSIDL_FLAG_DONT_VERIFY 0x4000
#define CSIDL_FLAG_NO_ALIAS 0x1000
#define CSIDL_FLAG_PER_USER_INIT 0x0800
#define CSIDL_FLAG_MASK 0xFF00
#define SHCNE_RENAMEITEM 0x00000001L
#define SHCNE_CREATE 0x00000002L
#define SHCNE_DELETE 0x00000004L
#define SHCNE_MKDIR 0x00000008L
#define SHCNE_RMDIR 0x00000010L
#define SHCNE_MEDIAINSERTED 0x00000020L
#define SHCNE_MEDIAREMOVED 0x00000040L
#define SHCNE_DRIVEREMOVED 0x00000080L
#define SHCNE_DRIVEADD 0x00000100L
#define SHCNE_NETSHARE 0x00000200L
#define SHCNE_NETUNSHARE 0x00000400L
#define SHCNE_ATTRIBUTES 0x00000800L
#define SHCNE_UPDATEDIR 0x00001000L
#define SHCNE_UPDATEITEM 0x00002000L
#define SHCNE_SERVERDISCONNECT 0x00004000L
#define SHCNE_UPDATEIMAGE 0x00008000L
#define SHCNE_DRIVEADDGUI 0x00010000L
#define SHCNE_RENAMEFOLDER 0x00020000L
#define SHCNE_FREESPACE 0x00040000L
#define SHCNE_EXTENDED_EVENT 0x04000000L
#define SHCNE_ASSOCCHANGED 0x08000000L
#define SHCNE_DISKEVENTS 0x0002381FL
#define SHCNE_GLOBALEVENTS 0x0C0581E0L
#define SHCNE_ALLEVENTS 0x7FFFFFFFL
#define SHCNE_INTERRUPT 0x80000000L
#define SHCNEE_ORDERCHANGED 2L
#define SHCNEE_MSI_CHANGE 4L
#define SHCNEE_MSI_UNINSTALL 5L
#define SHCNF_IDLIST 0x0000
#define SHCNF_PATHA 0x0001
#define SHCNF_PRINTERA 0x0002
#define SHCNF_DWORD 0x0003
#define SHCNF_PATHW 0x0005
#define SHCNF_PRINTERW 0x0006
#define SHCNF_TYPE 0x00FF
#define SHCNF_FLUSH 0x1000
#define SHCNF_FLUSHNOWAIT 0x2000
#define SHCNF_PATH SHCNF_PATHA
#define SHCNF_PRINTER SHCNF_PRINTERA
#define SQL_NULL_DATA (-1)
#define SQL_DATA_AT_EXEC (-2)
#define SQL_SUCCESS 0
#define SQL_SUCCESS_WITH_INFO 1
#define SQL_NO_DATA 100
#define SQL_ERROR (-1)
#define SQL_INVALID_HANDLE (-2)
#define SQL_STILL_EXECUTING 2
#define SQL_NEED_DATA 99
#define SQL_NTS (-3)
#define SQL_NTSL (-3L)
#define SQL_MAX_MESSAGE_LENGTH 512
#define SQL_DATE_LEN 10
#define SQL_TIME_LEN 8 
#define SQL_TIMESTAMP_LEN 19 
#define SQL_HANDLE_ENV 1
#define SQL_HANDLE_DBC 2
#define SQL_HANDLE_STMT 3
#define SQL_HANDLE_DESC 4
#define SQL_ATTR_OUTPUT_NTS 10001
#define SQL_ATTR_AUTO_IPD 10001
#define SQL_ATTR_METADATA_ID 10014
#define SQL_ATTR_APP_ROW_DESC 10010
#define SQL_ATTR_APP_PARAM_DESC 10011
#define SQL_ATTR_IMP_ROW_DESC 10012
#define SQL_ATTR_IMP_PARAM_DESC 10013
#define SQL_ATTR_CURSOR_SCROLLABLE (-1)
#define SQL_ATTR_CURSOR_SENSITIVITY (-2)
#define SQL_NONSCROLLABLE 0
#define SQL_SCROLLABLE 1
#define SQL_DESC_COUNT 1001
#define SQL_DESC_TYPE 1002
#define SQL_DESC_LENGTH 1003
#define SQL_DESC_OCTET_LENGTH_PTR 1004
#define SQL_DESC_PRECISION 1005
#define SQL_DESC_SCALE 1006
#define SQL_DESC_DATETIME_INTERVAL_CODE 1007
#define SQL_DESC_NULLABLE 1008
#define SQL_DESC_INDICATOR_PTR 1009
#define SQL_DESC_DATA_PTR 1010
#define SQL_DESC_NAME 1011
#define SQL_DESC_UNNAMED 1012
#define SQL_DESC_OCTET_LENGTH 1013
#define SQL_DESC_ALLOC_TYPE 1099
#define SQL_DIAG_RETURNCODE 1
#define SQL_DIAG_NUMBER 2
#define SQL_DIAG_ROW_COUNT 3
#define SQL_DIAG_SQLSTATE 4
#define SQL_DIAG_NATIVE 5
#define SQL_DIAG_MESSAGE_TEXT 6
#define SQL_DIAG_DYNAMIC_FUNCTION 7
#define SQL_DIAG_CLASS_ORIGIN 8
#define SQL_DIAG_SUBCLASS_ORIGIN 9
#define SQL_DIAG_CONNECTION_NAME 10
#define SQL_DIAG_SERVER_NAME 11
#define SQL_DIAG_DYNAMIC_FUNCTION_CODE 12
#define SQL_DIAG_ALTER_DOMAIN 3
#define SQL_DIAG_ALTER_TABLE 4
#define SQL_DIAG_CALL 7
#define SQL_DIAG_CREATE_ASSERTION 6
#define SQL_DIAG_CREATE_CHARACTER_SET 8
#define SQL_DIAG_CREATE_COLLATION 10
#define SQL_DIAG_CREATE_DOMAIN 23
#define SQL_DIAG_CREATE_INDEX (-1)
#define SQL_DIAG_CREATE_SCHEMA 64
#define SQL_DIAG_CREATE_TABLE 77
#define SQL_DIAG_CREATE_TRANSLATION 79
#define SQL_DIAG_CREATE_VIEW 84
#define SQL_DIAG_DELETE_WHERE 19
#define SQL_DIAG_DROP_ASSERTION 24
#define SQL_DIAG_DROP_CHARACTER_SET 25
#define SQL_DIAG_DROP_COLLATION 26
#define SQL_DIAG_DROP_DOMAIN 27
#define SQL_DIAG_DROP_INDEX (-2)
#define SQL_DIAG_DROP_SCHEMA 31
#define SQL_DIAG_DROP_TABLE 32
#define SQL_DIAG_DROP_TRANSLATION 33
#define SQL_DIAG_DROP_VIEW 36
#define SQL_DIAG_DYNAMIC_DELETE_CURSOR 38
#define SQL_DIAG_DYNAMIC_UPDATE_CURSOR 81
#define SQL_DIAG_GRANT 48
#define SQL_DIAG_INSERT 50
#define SQL_DIAG_REVOKE 59
#define SQL_DIAG_SELECT_CURSOR 85
#define SQL_DIAG_UNKNOWN_STATEMENT 0
#define SQL_DIAG_UPDATE_WHERE 82
#define SQL_UNKNOWN_TYPE 0
#define SQL_CHAR 1
#define SQL_NUMERIC 2
#define SQL_DECIMAL 3
#define SQL_INTEGER 4
#define SQL_SMALLINT 5
#define SQL_FLOAT 6
#define SQL_REAL 7
#define SQL_DOUBLE 8
#define SQL_DATETIME 9
#define SQL_VARCHAR 12
#define SQL_TYPE_DATE 91
#define SQL_TYPE_TIME 92
#define SQL_TYPE_TIMESTAMP 93
#define SQL_UNSPECIFIED 0
#define SQL_INSENSITIVE 1
#define SQL_SENSITIVE 2
#define SQL_ALL_TYPES 0
#define SQL_DEFAULT 99
#define SQL_ARD_TYPE (-99)
#define SQL_CODE_DATE 1
#define SQL_CODE_TIME 2
#define SQL_CODE_TIMESTAMP 3
#define SQL_FALSE 0
#define SQL_TRUE 1
#define SQL_NO_NULLS 0
#define SQL_NULLABLE 1
#define SQL_NULLABLE_UNKNOWN 2
#define SQL_PRED_NONE 0
#define SQL_PRED_CHAR 1
#define SQL_PRED_BASIC 2
#define SQL_NAMED 0
#define SQL_UNNAMED 1
#define SQL_DESC_ALLOC_AUTO 1
#define SQL_DESC_ALLOC_USER 2
#define SQL_CLOSE 0
#define SQL_DROP 1
#define SQL_UNBIND 2
#define SQL_RESET_PARAMS 3
#define SQL_FETCH_NEXT 1
#define SQL_FETCH_FIRST 2
#define SQL_FETCH_LAST 3
#define SQL_FETCH_PRIOR 4
#define SQL_FETCH_ABSOLUTE 5
#define SQL_FETCH_RELATIVE 6
#define SQL_COMMIT 0
#define SQL_ROLLBACK 1
#define SQL_NULL_HENV NULL_PTR
#define SQL_NULL_HDBC NULL_PTR
#define SQL_NULL_HSTMT NULL_PTR
#define SQL_NULL_HDESC NULL_PTR
#define SQL_NULL_HANDLE NULL_PTR
#define SQL_SCOPE_CURROW 0
#define SQL_SCOPE_TRANSACTION 1
#define SQL_SCOPE_SESSION 2
#define SQL_PC_UNKNOWN 0
#define SQL_PC_NON_PSEUDO 1
#define SQL_PC_PSEUDO 2
#define SQL_ROW_IDENTIFIER 1
#define SQL_INDEX_UNIQUE 0
#define SQL_INDEX_ALL 1
#define SQL_INDEX_CLUSTERED 1
#define SQL_INDEX_HASHED 2
#define SQL_INDEX_OTHER 3
#define SQL_API_SQLALLOCCONNECT 1
#define SQL_API_SQLALLOCENV 2
#define SQL_API_SQLALLOCHANDLE 1001
#define SQL_API_SQLALLOCSTMT 3
#define SQL_API_SQLBINDCOL 4
#define SQL_API_SQLBINDPARAM 1002
#define SQL_API_SQLCANCEL 5
#define SQL_API_SQLCLOSECURSOR 1003
#define SQL_API_SQLCOLATTRIBUTE 6
#define SQL_API_SQLCOLUMNS 40
#define SQL_API_SQLCONNECT 7
#define SQL_API_SQLCOPYDESC 1004
#define SQL_API_SQLDATASOURCES 57
#define SQL_API_SQLDESCRIBECOL 8
#define SQL_API_SQLDISCONNECT 9
#define SQL_API_SQLENDTRAN 1005
#define SQL_API_SQLERROR 10
#define SQL_API_SQLEXECDIRECT 11
#define SQL_API_SQLEXECUTE 12
#define SQL_API_SQLFETCH 13
#define SQL_API_SQLFETCHSCROLL 1021
#define SQL_API_SQLFREECONNECT 14
#define SQL_API_SQLFREEENV 15
#define SQL_API_SQLFREEHANDLE 1006
#define SQL_API_SQLFREESTMT 16
#define SQL_API_SQLGETCONNECTATTR 1007
#define SQL_API_SQLGETCONNECTOPTION 42
#define SQL_API_SQLGETCURSORNAME 17
#define SQL_API_SQLGETDATA 43
#define SQL_API_SQLGETDESCFIELD 1008
#define SQL_API_SQLGETDESCREC 1009
#define SQL_API_SQLGETDIAGFIELD 1010
#define SQL_API_SQLGETDIAGREC 1011
#define SQL_API_SQLGETENVATTR 1012
#define SQL_API_SQLGETFUNCTIONS 44
#define SQL_API_SQLGETINFO 45
#define SQL_API_SQLGETSTMTATTR 1014
#define SQL_API_SQLGETSTMTOPTION 46
#define SQL_API_SQLGETTYPEINFO 47
#define SQL_API_SQLNUMRESULTCOLS 18
#define SQL_API_SQLPARAMDATA 48
#define SQL_API_SQLPREPARE 19
#define SQL_API_SQLPUTDATA 49
#define SQL_API_SQLROWCOUNT 20
#define SQL_API_SQLSETCONNECTATTR 1016
#define SQL_API_SQLSETCONNECTOPTION 50
#define SQL_API_SQLSETCURSORNAME 21
#define SQL_API_SQLSETDESCFIELD 1017
#define SQL_API_SQLSETDESCREC 1018
#define SQL_API_SQLSETENVATTR 1019
#define SQL_API_SQLSETPARAM 22
#define SQL_API_SQLSETSTMTATTR 1020
#define SQL_API_SQLSETSTMTOPTION 51
#define SQL_API_SQLSPECIALCOLUMNS 52
#define SQL_API_SQLSTATISTICS 53
#define SQL_API_SQLTABLES 54
#define SQL_API_SQLTRANSACT 23
#define SQL_MAX_DRIVER_CONNECTIONS 0
#define SQL_MAXIMUM_DRIVER_CONNECTIONS SQL_MAX_DRIVER_CONNECTIONS
#define SQL_MAX_CONCURRENT_ACTIVITIES 1
#define SQL_MAXIMUM_CONCURRENT_ACTIVITIES SQL_MAX_CONCURRENT_ACTIVITIES
#define SQL_DATA_SOURCE_NAME 2
#define SQL_FETCH_DIRECTION 8
#define SQL_SERVER_NAME 13
#define SQL_SEARCH_PATTERN_ESCAPE 14
#define SQL_DBMS_NAME 17
#define SQL_DBMS_VER 18
#define SQL_ACCESSIBLE_TABLES 19
#define SQL_ACCESSIBLE_PROCEDURES 20
#define SQL_CURSOR_COMMIT_BEHAVIOR 23
#define SQL_DATA_SOURCE_READ_ONLY 25
#define SQL_DEFAULT_TXN_ISOLATION 26
#define SQL_IDENTIFIER_CASE 28
#define SQL_IDENTIFIER_QUOTE_CHAR 29
#define SQL_MAX_COLUMN_NAME_LEN 30
#define SQL_MAXIMUM_COLUMN_NAME_LENGTH SQL_MAX_COLUMN_NAME_LEN
#define SQL_MAX_CURSOR_NAME_LEN 31
#define SQL_MAXIMUM_CURSOR_NAME_LENGTH SQL_MAX_CURSOR_NAME_LEN
#define SQL_MAX_SCHEMA_NAME_LEN 32
#define SQL_MAXIMUM_SCHEMA_NAME_LENGTH SQL_MAX_SCHEMA_NAME_LEN
#define SQL_MAX_CATALOG_NAME_LEN 34
#define SQL_MAXIMUM_CATALOG_NAME_LENGTH SQL_MAX_CATALOG_NAME_LEN
#define SQL_MAX_TABLE_NAME_LEN 35
#define SQL_SCROLL_CONCURRENCY 43
#define SQL_TXN_CAPABLE 46
#define SQL_TRANSACTION_CAPABLE SQL_TXN_CAPABLE
#define SQL_USER_NAME 47
#define SQL_TXN_ISOLATION_OPTION 72
#define SQL_TRANSACTION_ISOLATION_OPTION SQL_TXN_ISOLATION_OPTION
#define SQL_INTEGRITY 73
#define SQL_GETDATA_EXTENSIONS 81
#define SQL_NULL_COLLATION 85
#define SQL_ALTER_TABLE 86
#define SQL_ORDER_BY_COLUMNS_IN_SELECT 90
#define SQL_SPECIAL_CHARACTERS 94
#define SQL_MAX_COLUMNS_IN_GROUP_BY 97
#define SQL_MAXIMUM_COLUMNS_IN_GROUP_BY SQL_MAX_COLUMNS_IN_GROUP_BY
#define SQL_MAX_COLUMNS_IN_INDEX 98
#define SQL_MAXIMUM_COLUMNS_IN_INDEX SQL_MAX_COLUMNS_IN_INDEX
#define SQL_MAX_COLUMNS_IN_ORDER_BY 99
#define SQL_MAXIMUM_COLUMNS_IN_ORDER_BY SQL_MAX_COLUMNS_IN_ORDER_BY
#define SQL_MAX_COLUMNS_IN_SELECT 100
#define SQL_MAXIMUM_COLUMNS_IN_SELECT SQL_MAX_COLUMNS_IN_SELECT
#define SQL_MAX_COLUMNS_IN_TABLE 101
#define SQL_MAX_INDEX_SIZE 102
#define SQL_MAXIMUM_INDEX_SIZE SQL_MAX_INDEX_SIZE
#define SQL_MAX_ROW_SIZE 104
#define SQL_MAXIMUM_ROW_SIZE SQL_MAX_ROW_SIZE
#define SQL_MAX_STATEMENT_LEN 105
#define SQL_MAXIMUM_STATEMENT_LENGTH SQL_MAX_STATEMENT_LEN
#define SQL_MAX_TABLES_IN_SELECT 106
#define SQL_MAXIMUM_TABLES_IN_SELECT SQL_MAX_TABLES_IN_SELECT
#define SQL_MAX_USER_NAME_LEN 107
#define SQL_MAXIMUM_USER_NAME_LENGTH SQL_MAX_USER_NAME_LEN
#define SQL_OJ_CAPABILITIES 115
#define SQL_OUTER_JOIN_CAPABILITIES SQL_OJ_CAPABILITIES
#define SQL_XOPEN_CLI_YEAR 10000
#define SQL_CURSOR_SENSITIVITY 10001
#define SQL_DESCRIBE_PARAMETER 10002
#define SQL_CATALOG_NAME 10003
#define SQL_COLLATION_SEQ 10004
#define SQL_MAX_IDENTIFIER_LEN 10005
#define SQL_MAXIMUM_IDENTIFIER_LENGTH SQL_MAX_IDENTIFIER_LEN
#define SQL_AT_ADD_COLUMN 0x00000001L
#define SQL_AT_DROP_COLUMN 0x00000002L
#define SQL_AT_ADD_CONSTRAINT 0x00000008L
#define SQL_AM_NONE 0
#define SQL_AM_CONNECTION 1
#define SQL_AM_STATEMENT 2
#define SQL_CB_DELETE 0
#define SQL_CB_CLOSE 1
#define SQL_CB_PRESERVE 2
#define SQL_FD_FETCH_NEXT 0x00000001L
#define SQL_FD_FETCH_FIRST 0x00000002L
#define SQL_FD_FETCH_LAST 0x00000004L
#define SQL_FD_FETCH_PRIOR 0x00000008L
#define SQL_FD_FETCH_ABSOLUTE 0x00000010L
#define SQL_FD_FETCH_RELATIVE 0x00000020L
#define SQL_GD_ANY_COLUMN 0x00000001L
#define SQL_GD_ANY_ORDER 0x00000002L
#define SQL_IC_UPPER 1
#define SQL_IC_LOWER 2
#define SQL_IC_SENSITIVE 3
#define SQL_IC_MIXED 4
#define SQL_OJ_LEFT 0x00000001L
#define SQL_OJ_RIGHT 0x00000002L
#define SQL_OJ_FULL 0x00000004L
#define SQL_OJ_NESTED 0x00000008L
#define SQL_OJ_NOT_ORDERED 0x00000010L
#define SQL_OJ_INNER 0x00000020L
#define SQL_OJ_ALL_COMPARISON_OPS 0x00000040L
#define SQL_SCCO_READ_ONLY 0x00000001L
#define SQL_SCCO_LOCK 0x00000002L
#define SQL_SCCO_OPT_ROWVER 0x00000004L
#define SQL_SCCO_OPT_VALUES 0x00000008L
#define SQL_TC_NONE 0
#define SQL_TC_DML 1
#define SQL_TC_ALL 2
#define SQL_TC_DDL_COMMIT 3
#define SQL_TC_DDL_IGNORE 4
#define SQL_TXN_READ_UNCOMMITTED 0x00000001L
#define SQL_TRANSACTION_READ_UNCOMMITTED SQL_TXN_READ_UNCOMMITTED
#define SQL_TXN_READ_COMMITTED 0x00000002L
#define SQL_TRANSACTION_READ_COMMITTED SQL_TXN_READ_COMMITTED
#define SQL_TXN_REPEATABLE_READ 0x00000004L
#define SQL_TRANSACTION_REPEATABLE_READ SQL_TXN_REPEATABLE_READ
#define SQL_TXN_SERIALIZABLE 0x00000008L
#define SQL_TRANSACTION_SERIALIZABLE SQL_TXN_SERIALIZABLE
#define SQL_NC_HIGH 0
#define SQL_NC_LOW 1
#define SQL_SPEC_MAJOR 3 
#define SQL_SPEC_MINOR 52 
#define SQL_SPEC_STRING "03.52" 
#define SQL_SQLSTATE_SIZE 5 
#define SQL_MAX_DSN_LENGTH 32 
#define SQL_MAX_OPTION_STRING_LENGTH 256
#define SQL_NO_DATA_FOUND SQL_NO_DATA
#define SQL_HANDLE_SENV 5
#define SQL_ATTR_ODBC_VERSION 200
#define SQL_ATTR_CONNECTION_POOLING 201
#define SQL_ATTR_CP_MATCH 202
#define SQL_CP_OFF 0U
#define SQL_CP_ONE_PER_DRIVER 1U
#define SQL_CP_ONE_PER_HENV 2U
#define SQL_CP_DEFAULT SQL_CP_OFF
#define SQL_CP_STRICT_MATCH 0U
#define SQL_CP_RELAXED_MATCH 1U
#define SQL_CP_MATCH_DEFAULT SQL_CP_STRICT_MATCH
#define SQL_OV_ODBC2 2U
#define SQL_OV_ODBC3 3U
#define SQL_ACCESS_MODE 101
#define SQL_AUTOCOMMIT 102
#define SQL_LOGIN_TIMEOUT 103
#define SQL_OPT_TRACE 104
#define SQL_OPT_TRACEFILE 105
#define SQL_TRANSLATE_DLL 106
#define SQL_TRANSLATE_OPTION 107
#define SQL_TXN_ISOLATION 108
#define SQL_CURRENT_QUALIFIER 109
#define SQL_ODBC_CURSORS 110
#define SQL_QUIET_MODE 111
#define SQL_PACKET_SIZE 112
#define SQL_ATTR_ACCESS_MODE SQL_ACCESS_MODE
#define SQL_ATTR_AUTOCOMMIT SQL_AUTOCOMMIT
#define SQL_ATTR_CONNECTION_TIMEOUT 113
#define SQL_ATTR_CURRENT_CATALOG SQL_CURRENT_QUALIFIER
#define SQL_ATTR_DISCONNECT_BEHAVIOR 114
#define SQL_ATTR_ENLIST_IN_DTC 1207
#define SQL_ATTR_ENLIST_IN_XA 1208
#define SQL_ATTR_LOGIN_TIMEOUT SQL_LOGIN_TIMEOUT
#define SQL_ATTR_ODBC_CURSORS SQL_ODBC_CURSORS
#define SQL_ATTR_PACKET_SIZE SQL_PACKET_SIZE
#define SQL_ATTR_QUIET_MODE SQL_QUIET_MODE
#define SQL_ATTR_TRACE SQL_OPT_TRACE
#define SQL_ATTR_TRACEFILE SQL_OPT_TRACEFILE
#define SQL_ATTR_TRANSLATE_LIB SQL_TRANSLATE_DLL
#define SQL_ATTR_TRANSLATE_OPTION SQL_TRANSLATE_OPTION
#define SQL_ATTR_TXN_ISOLATION SQL_TXN_ISOLATION
#define SQL_ATTR_CONNECTION_DEAD 1209 
#define SQL_MODE_READ_WRITE 0U
#define SQL_MODE_READ_ONLY 1U
#define SQL_MODE_DEFAULT SQL_MODE_READ_WRITE
#define SQL_AUTOCOMMIT_OFF 0U
#define SQL_AUTOCOMMIT_ON 1U
#define SQL_AUTOCOMMIT_DEFAULT SQL_AUTOCOMMIT_ON
#define SQL_LOGIN_TIMEOUT_DEFAULT 15U
#define SQL_OPT_TRACE_OFF 0U
#define SQL_OPT_TRACE_ON 1U
#define SQL_OPT_TRACE_DEFAULT SQL_OPT_TRACE_OFF
#define SQL_OPT_TRACE_FILE_DEFAULT "\\SQL.LOG"
#define SQL_CUR_USE_IF_NEEDED 0U
#define SQL_CUR_USE_ODBC 1U
#define SQL_CUR_USE_DRIVER 2U
#define SQL_CUR_DEFAULT SQL_CUR_USE_DRIVER
#define SQL_DB_RETURN_TO_POOL 0U
#define SQL_DB_DISCONNECT 1U
#define SQL_DB_DEFAULT SQL_DB_RETURN_TO_POOL
#define SQL_DTC_DONE 0L
#define SQL_CD_TRUE 1L 
#define SQL_CD_FALSE 0L 
#define SQL_QUERY_TIMEOUT 0
#define SQL_MAX_ROWS 1
#define SQL_NOSCAN 2
#define SQL_MAX_LENGTH 3
#define SQL_ASYNC_ENABLE 4 
#define SQL_BIND_TYPE 5
#define SQL_CURSOR_TYPE 6
#define SQL_CONCURRENCY 7
#define SQL_KEYSET_SIZE 8
#define SQL_ROWSET_SIZE 9
#define SQL_SIMULATE_CURSOR 10
#define SQL_RETRIEVE_DATA 11
#define SQL_USE_BOOKMARKS 12
#define SQL_GET_BOOKMARK 13 
#define SQL_ROW_NUMBER 14 
#define SQL_ATTR_ASYNC_ENABLE 4
#define SQL_ATTR_CONCURRENCY SQL_CONCURRENCY
#define SQL_ATTR_CURSOR_TYPE SQL_CURSOR_TYPE
#define SQL_ATTR_ENABLE_AUTO_IPD 15
#define SQL_ATTR_FETCH_BOOKMARK_PTR 16
#define SQL_ATTR_KEYSET_SIZE SQL_KEYSET_SIZE
#define SQL_ATTR_MAX_LENGTH SQL_MAX_LENGTH
#define SQL_ATTR_MAX_ROWS SQL_MAX_ROWS
#define SQL_ATTR_NOSCAN SQL_NOSCAN
#define SQL_ATTR_PARAM_BIND_OFFSET_PTR 17
#define SQL_ATTR_PARAM_BIND_TYPE 18
#define SQL_ATTR_PARAM_OPERATION_PTR 19
#define SQL_ATTR_PARAM_STATUS_PTR 20
#define SQL_ATTR_PARAMS_PROCESSED_PTR 21
#define SQL_ATTR_PARAMSET_SIZE 22
#define SQL_ATTR_QUERY_TIMEOUT SQL_QUERY_TIMEOUT
#define SQL_ATTR_RETRIEVE_DATA SQL_RETRIEVE_DATA
#define SQL_ATTR_ROW_BIND_OFFSET_PTR 23
#define SQL_ATTR_ROW_BIND_TYPE SQL_BIND_TYPE
#define SQL_ATTR_ROW_NUMBER SQL_ROW_NUMBER 
#define SQL_ATTR_ROW_OPERATION_PTR 24
#define SQL_ATTR_ROW_STATUS_PTR 25
#define SQL_ATTR_ROWS_FETCHED_PTR 26
#define SQL_ATTR_ROW_ARRAY_SIZE 27
#define SQL_ATTR_SIMULATE_CURSOR SQL_SIMULATE_CURSOR
#define SQL_ATTR_USE_BOOKMARKS SQL_USE_BOOKMARKS
#define SQL_LIKE_ONLY 1
#define SQL_COL_PRED_CHAR SQL_LIKE_ONLY
#define SQL_ALL_EXCEPT_LIKE 2
#define SQL_COL_PRED_BASIC SQL_ALL_EXCEPT_LIKE
#define SQL_IS_POINTER (-4)
#define SQL_IS_UINTEGER (-5)
#define SQL_IS_INTEGER (-6)
#define SQL_IS_USMALLINT (-7)
#define SQL_IS_SMALLINT (-8)
#define SQL_PARAM_BIND_BY_COLUMN 0U
#define SQL_PARAM_BIND_TYPE_DEFAULT SQL_PARAM_BIND_BY_COLUMN
#define SQL_QUERY_TIMEOUT_DEFAULT 0U
#define SQL_MAX_ROWS_DEFAULT 0U
#define SQL_NOSCAN_OFF 0U 
#define SQL_NOSCAN_ON 1U 
#define SQL_NOSCAN_DEFAULT SQL_NOSCAN_OFF
#define SQL_MAX_LENGTH_DEFAULT 0U
#define SQL_ASYNC_ENABLE_OFF 0U
#define SQL_ASYNC_ENABLE_ON 1U
#define SQL_ASYNC_ENABLE_DEFAULT SQL_ASYNC_ENABLE_OFF
#define SQL_BIND_BY_COLUMN 0U
#define SQL_BIND_TYPE_DEFAULT SQL_BIND_BY_COLUMN 
#define SQL_CONCUR_READ_ONLY 1
#define SQL_CONCUR_LOCK 2
#define SQL_CONCUR_ROWVER 3
#define SQL_CONCUR_VALUES 4
#define SQL_CONCUR_DEFAULT SQL_CONCUR_READ_ONLY 
#define SQL_CURSOR_FORWARD_ONLY 0U
#define SQL_CURSOR_KEYSET_DRIVEN 1U
#define SQL_CURSOR_DYNAMIC 2U
#define SQL_CURSOR_STATIC 3U
#define SQL_CURSOR_TYPE_DEFAULT SQL_CURSOR_FORWARD_ONLY 
#define SQL_ROWSET_SIZE_DEFAULT 1U
#define SQL_KEYSET_SIZE_DEFAULT 0U
#define SQL_SC_NON_UNIQUE 0U
#define SQL_SC_TRY_UNIQUE 1U
#define SQL_SC_UNIQUE 2U
#define SQL_RD_OFF 0U
#define SQL_RD_ON 1U
#define SQL_RD_DEFAULT SQL_RD_ON
#define SQL_UB_OFF 0U
#define SQL_UB_ON 01U
#define SQL_UB_DEFAULT SQL_UB_OFF
#define SQL_UB_FIXED SQL_UB_ON
#define SQL_UB_VARIABLE 2U
#define SQL_DESC_ARRAY_SIZE 20
#define SQL_DESC_ARRAY_STATUS_PTR 21
#define SQL_COLUMN_AUTO_INCREMENT 11
#define SQL_DESC_AUTO_UNIQUE_VALUE SQL_COLUMN_AUTO_INCREMENT
#define SQL_DESC_BASE_COLUMN_NAME 22
#define SQL_DESC_BASE_TABLE_NAME 23
#define SQL_DESC_BIND_OFFSET_PTR 24
#define SQL_DESC_BIND_TYPE 25
#define SQL_COLUMN_CASE_SENSITIVE 12
#define SQL_DESC_CASE_SENSITIVE SQL_COLUMN_CASE_SENSITIVE
#define SQL_COLUMN_QUALIFIER_NAME 17
#define SQL_DESC_CATALOG_NAME SQL_COLUMN_QUALIFIER_NAME
#define SQL_COLUMN_TYPE 2
#define SQL_DESC_CONCISE_TYPE SQL_COLUMN_TYPE
#define SQL_DESC_DATETIME_INTERVAL_PRECISION 26
#define SQL_COLUMN_DISPLAY_SIZE 6
#define SQL_DESC_DISPLAY_SIZE SQL_COLUMN_DISPLAY_SIZE
#define SQL_COLUMN_MONEY 9
#define SQL_DESC_FIXED_PREC_SCALE SQL_COLUMN_MONEY
#define SQL_COLUMN_LABEL 18
#define SQL_DESC_LABEL SQL_COLUMN_LABEL
#define SQL_DESC_LITERAL_PREFIX 27
#define SQL_DESC_LITERAL_SUFFIX 28
#define SQL_DESC_LOCAL_TYPE_NAME 29
#define SQL_DESC_MAXIMUM_SCALE 30
#define SQL_DESC_MINIMUM_SCALE 31
#define SQL_DESC_NUM_PREC_RADIX 32
#define SQL_DESC_PARAMETER_TYPE 33
#define SQL_DESC_ROWS_PROCESSED_PTR 34
#define SQL_DESC_ROWVER 35
#define SQL_COLUMN_OWNER_NAME 16
#define SQL_DESC_SCHEMA_NAME SQL_COLUMN_OWNER_NAME
#define SQL_COLUMN_SEARCHABLE 13
#define SQL_DESC_SEARCHABLE SQL_COLUMN_SEARCHABLE
#define SQL_COLUMN_TYPE_NAME 14
#define SQL_DESC_TYPE_NAME SQL_COLUMN_TYPE_NAME
#define SQL_COLUMN_TABLE_NAME 15
#define SQL_DESC_TABLE_NAME SQL_COLUMN_TABLE_NAME
#define SQL_COLUMN_UNSIGNED 8
#define SQL_DESC_UNSIGNED SQL_COLUMN_UNSIGNED
#define SQL_COLUMN_UPDATABLE 10
#define SQL_DESC_UPDATABLE SQL_COLUMN_UPDATABLE
#define SQL_DIAG_CURSOR_ROW_COUNT (-1249)
#define SQL_DIAG_ROW_NUMBER (-1248)
#define SQL_DIAG_COLUMN_NUMBER (-1247)
#define SQL_DATE 9
#define SQL_INTERVAL 10
#define SQL_TIME 10
#define SQL_TIMESTAMP 11
#define SQL_LONGVARCHAR (-1)
#define SQL_BINARY (-2)
#define SQL_VARBINARY (-3)
#define SQL_LONGVARBINARY (-4)
#define SQL_BIGINT (-5)
#define SQL_TINYINT (-6)
#define SQL_BIT (-7)
#define SQL_GUID (-11)
#define SQL_CODE_YEAR 1
#define SQL_CODE_MONTH 2
#define SQL_CODE_DAY 3
#define SQL_CODE_HOUR 4
#define SQL_CODE_MINUTE 5
#define SQL_CODE_SECOND 6
#define SQL_CODE_YEAR_TO_MONTH 7
#define SQL_CODE_DAY_TO_HOUR 8
#define SQL_CODE_DAY_TO_MINUTE 9
#define SQL_CODE_DAY_TO_SECOND 10
#define SQL_CODE_HOUR_TO_MINUTE 11
#define SQL_CODE_HOUR_TO_SECOND 12
#define SQL_CODE_MINUTE_TO_SECOND 13
#define SQL_INTERVAL_YEAR (100 + SQL_CODE_YEAR)
#define SQL_INTERVAL_MONTH (100 + SQL_CODE_MONTH)
#define SQL_INTERVAL_DAY (100 + SQL_CODE_DAY)
#define SQL_INTERVAL_HOUR (100 + SQL_CODE_HOUR)
#define SQL_INTERVAL_MINUTE (100 + SQL_CODE_MINUTE)
#define SQL_INTERVAL_SECOND (100 + SQL_CODE_SECOND)
#define SQL_INTERVAL_YEAR_TO_MONTH (100 + SQL_CODE_YEAR_TO_MONTH)
#define SQL_INTERVAL_DAY_TO_HOUR (100 + SQL_CODE_DAY_TO_HOUR)
#define SQL_INTERVAL_DAY_TO_MINUTE (100 + SQL_CODE_DAY_TO_MINUTE)
#define SQL_INTERVAL_DAY_TO_SECOND (100 + SQL_CODE_DAY_TO_SECOND)
#define SQL_INTERVAL_HOUR_TO_MINUTE (100 + SQL_CODE_HOUR_TO_MINUTE)
#define SQL_INTERVAL_HOUR_TO_SECOND (100 + SQL_CODE_HOUR_TO_SECOND)
#define SQL_INTERVAL_MINUTE_TO_SECOND (100 + SQL_CODE_MINUTE_TO_SECOND)
#define SQL_WCHAR (-8)
#define SQL_UNICODE SQL_WCHAR
#define SQL_WVARCHAR (-9)
#define SQL_UNICODE_VARCHAR SQL_WVARCHAR
#define SQL_WLONGVARCHAR (-10)
#define SQL_UNICODE_LONGVARCHAR SQL_WLONGVARCHAR
#define SQL_UNICODE_CHAR SQL_WCHAR
#define SQL_C_CHAR SQL_CHAR 
#define SQL_C_LONG SQL_INTEGER 
#define SQL_C_SHORT SQL_SMALLINT 
#define SQL_C_FLOAT SQL_REAL 
#define SQL_C_DOUBLE SQL_DOUBLE 
#define SQL_C_NUMERIC SQL_NUMERIC
#define SQL_C_DEFAULT 99
#define SQL_SIGNED_OFFSET (-20)
#define SQL_UNSIGNED_OFFSET (-22)
#define SQL_C_DATE SQL_DATE
#define SQL_C_TIME SQL_TIME
#define SQL_C_TIMESTAMP SQL_TIMESTAMP
#define SQL_C_TYPE_DATE SQL_TYPE_DATE
#define SQL_C_TYPE_TIME SQL_TYPE_TIME
#define SQL_C_TYPE_TIMESTAMP SQL_TYPE_TIMESTAMP
#define SQL_C_INTERVAL_YEAR SQL_INTERVAL_YEAR
#define SQL_C_INTERVAL_MONTH SQL_INTERVAL_MONTH
#define SQL_C_INTERVAL_DAY SQL_INTERVAL_DAY
#define SQL_C_INTERVAL_HOUR SQL_INTERVAL_HOUR
#define SQL_C_INTERVAL_MINUTE SQL_INTERVAL_MINUTE
#define SQL_C_INTERVAL_SECOND SQL_INTERVAL_SECOND
#define SQL_C_INTERVAL_YEAR_TO_MONTH SQL_INTERVAL_YEAR_TO_MONTH
#define SQL_C_INTERVAL_DAY_TO_HOUR SQL_INTERVAL_DAY_TO_HOUR
#define SQL_C_INTERVAL_DAY_TO_MINUTE SQL_INTERVAL_DAY_TO_MINUTE
#define SQL_C_INTERVAL_DAY_TO_SECOND SQL_INTERVAL_DAY_TO_SECOND
#define SQL_C_INTERVAL_HOUR_TO_MINUTE SQL_INTERVAL_HOUR_TO_MINUTE
#define SQL_C_INTERVAL_HOUR_TO_SECOND SQL_INTERVAL_HOUR_TO_SECOND
#define SQL_C_INTERVAL_MINUTE_TO_SECOND SQL_INTERVAL_MINUTE_TO_SECOND
#define SQL_C_BINARY SQL_BINARY
#define SQL_C_BIT SQL_BIT
#define SQL_C_SBIGINT (SQL_BIGINT+SQL_SIGNED_OFFSET) 
#define SQL_C_UBIGINT (SQL_BIGINT+SQL_UNSIGNED_OFFSET) 
#define SQL_C_TINYINT SQL_TINYINT
#define SQL_C_SLONG (SQL_C_LONG+SQL_SIGNED_OFFSET) 
#define SQL_C_SSHORT (SQL_C_SHORT+SQL_SIGNED_OFFSET) 
#define SQL_C_STINYINT (SQL_TINYINT+SQL_SIGNED_OFFSET) 
#define SQL_C_ULONG (SQL_C_LONG+SQL_UNSIGNED_OFFSET) 
#define SQL_C_USHORT (SQL_C_SHORT+SQL_UNSIGNED_OFFSET) 
#define SQL_C_UTINYINT (SQL_TINYINT+SQL_UNSIGNED_OFFSET) 
#define SQL_C_BOOKMARK SQL_C_ULONG 
#define SQL_C_GUID SQL_GUID
#define SQL_TYPE_NULL 0
#define SQL_C_VARBOOKMARK SQL_C_BINARY
#define SQL_NO_ROW_NUMBER (-1)
#define SQL_NO_COLUMN_NUMBER (-1)
#define SQL_ROW_NUMBER_UNKNOWN (-2)
#define SQL_COLUMN_NUMBER_UNKNOWN (-2)
#define SQL_DEFAULT_PARAM (-5)
#define SQL_IGNORE (-6)
#define SQL_COLUMN_IGNORE SQL_IGNORE
#define SQL_LEN_DATA_AT_EXEC_OFFSET (-100)
#define SQL_LEN_BINARY_ATTR_OFFSET (-100)
#define SQL_PARAM_INPUT_OUTPUT 2
#define SQL_PARAM_TYPE_DEFAULT SQL_PARAM_INPUT_OUTPUT
#define SQL_SETPARAM_VALUE_MAX (-1L)
#define SQL_COLUMN_COUNT 0
#define SQL_COLUMN_NAME 1
#define SQL_COLUMN_LENGTH 3
#define SQL_COLUMN_PRECISION 4
#define SQL_COLUMN_SCALE 5
#define SQL_COLUMN_NULLABLE 7
#define SQL_COLATT_OPT_MAX SQL_COLUMN_LABEL
#define SQL_COLATT_OPT_MIN SQL_COLUMN_COUNT
#define SQL_ATTR_READONLY 0
#define SQL_ATTR_WRITE 1
#define SQL_ATTR_READWRITE_UNKNOWN 2
#define SQL_UNSEARCHABLE 0
#define SQL_SEARCHABLE 3
#define SQL_PRED_SEARCHABLE SQL_SEARCHABLE
#define SQL_NO_TOTAL (-4)
#define SQL_API_SQLALLOCHANDLESTD 73
#define SQL_API_SQLBULKOPERATIONS 24
#define SQL_API_SQLBINDPARAMETER 72
#define SQL_API_SQLBROWSECONNECT 55
#define SQL_API_SQLCOLATTRIBUTES 6
#define SQL_API_SQLCOLUMNPRIVILEGES 56
#define SQL_API_SQLDESCRIBEPARAM 58
#define SQL_API_SQLDRIVERCONNECT 41
#define SQL_API_SQLDRIVERS 71
#define SQL_API_SQLEXTENDEDFETCH 59
#define SQL_API_SQLFOREIGNKEYS 60
#define SQL_API_SQLMORERESULTS 61
#define SQL_API_SQLNATIVESQL 62
#define SQL_API_SQLNUMPARAMS 63
#define SQL_API_SQLPARAMOPTIONS 64
#define SQL_API_SQLPRIMARYKEYS 65
#define SQL_API_SQLPROCEDURECOLUMNS 66
#define SQL_API_SQLPROCEDURES 67
#define SQL_API_SQLSETPOS 68
#define SQL_API_SQLSETSCROLLOPTIONS 69
#define SQL_API_SQLTABLEPRIVILEGES 70
#define SQL_API_ALL_FUNCTIONS 0 
#define SQL_API_LOADBYORDINAL 199 
#define SQL_API_ODBC3_ALL_FUNCTIONS 999
#define SQL_API_ODBC3_ALL_FUNCTIONS_SIZE 250 
#define SQL_INFO_FIRST 0
#define SQL_ACTIVE_CONNECTIONS 0 
#define SQL_ACTIVE_STATEMENTS 1 
#define SQL_DRIVER_HDBC 3
#define SQL_DRIVER_HENV 4
#define SQL_DRIVER_HSTMT 5
#define SQL_DRIVER_NAME 6
#define SQL_DRIVER_VER 7
#define SQL_ODBC_API_CONFORMANCE 9
#define SQL_ODBC_VER 10
#define SQL_ROW_UPDATES 11
#define SQL_ODBC_SAG_CLI_CONFORMANCE 12
#define SQL_ODBC_SQL_CONFORMANCE 15
#define SQL_PROCEDURES 21
#define SQL_CONCAT_NULL_BEHAVIOR 22
#define SQL_CURSOR_ROLLBACK_BEHAVIOR 24
#define SQL_EXPRESSIONS_IN_ORDERBY 27
#define SQL_MAX_OWNER_NAME_LEN 32 
#define SQL_MAX_PROCEDURE_NAME_LEN 33
#define SQL_MAX_QUALIFIER_NAME_LEN 34 
#define SQL_MULT_RESULT_SETS 36
#define SQL_MULTIPLE_ACTIVE_TXN 37
#define SQL_OUTER_JOINS 38
#define SQL_OWNER_TERM 39
#define SQL_PROCEDURE_TERM 40
#define SQL_QUALIFIER_NAME_SEPARATOR 41
#define SQL_QUALIFIER_TERM 42
#define SQL_SCROLL_OPTIONS 44
#define SQL_TABLE_TERM 45
#define SQL_CONVERT_FUNCTIONS 48
#define SQL_NUMERIC_FUNCTIONS 49
#define SQL_STRING_FUNCTIONS 50
#define SQL_SYSTEM_FUNCTIONS 51
#define SQL_TIMEDATE_FUNCTIONS 52
#define SQL_CONVERT_BIGINT 53
#define SQL_CONVERT_BINARY 54
#define SQL_CONVERT_BIT 55
#define SQL_CONVERT_CHAR 56
#define SQL_CONVERT_DATE 57
#define SQL_CONVERT_DECIMAL 58
#define SQL_CONVERT_DOUBLE 59
#define SQL_CONVERT_FLOAT 60
#define SQL_CONVERT_INTEGER 61
#define SQL_CONVERT_LONGVARCHAR 62
#define SQL_CONVERT_NUMERIC 63
#define SQL_CONVERT_REAL 64
#define SQL_CONVERT_SMALLINT 65
#define SQL_CONVERT_TIME 66
#define SQL_CONVERT_TIMESTAMP 67
#define SQL_CONVERT_TINYINT 68
#define SQL_CONVERT_VARBINARY 69
#define SQL_CONVERT_VARCHAR 70
#define SQL_CONVERT_LONGVARBINARY 71
#define SQL_ODBC_SQL_OPT_IEF 73 
#define SQL_CORRELATION_NAME 74
#define SQL_NON_NULLABLE_COLUMNS 75
#define SQL_DRIVER_HLIB 76
#define SQL_DRIVER_ODBC_VER 77
#define SQL_LOCK_TYPES 78
#define SQL_POS_OPERATIONS 79
#define SQL_POSITIONED_STATEMENTS 80
#define SQL_BOOKMARK_PERSISTENCE 82
#define SQL_STATIC_SENSITIVITY 83
#define SQL_FILE_USAGE 84
#define SQL_COLUMN_ALIAS 87
#define SQL_GROUP_BY 88
#define SQL_KEYWORDS 89
#define SQL_OWNER_USAGE 91
#define SQL_QUALIFIER_USAGE 92
#define SQL_QUOTED_IDENTIFIER_CASE 93
#define SQL_SUBQUERIES 95
#define SQL_UNION 96
#define SQL_MAX_ROW_SIZE_INCLUDES_LONG 103
#define SQL_MAX_CHAR_LITERAL_LEN 108
#define SQL_TIMEDATE_ADD_INTERVALS 109
#define SQL_TIMEDATE_DIFF_INTERVALS 110
#define SQL_NEED_LONG_DATA_LEN 111
#define SQL_MAX_BINARY_LITERAL_LEN 112
#define SQL_LIKE_ESCAPE_CLAUSE 113
#define SQL_QUALIFIER_LOCATION 114
#define SQL_ACTIVE_ENVIRONMENTS 116
#define SQL_ALTER_DOMAIN 117
#define SQL_SQL_CONFORMANCE 118
#define SQL_DATETIME_LITERALS 119
#define SQL_ASYNC_MODE 10021 
#define SQL_BATCH_ROW_COUNT 120
#define SQL_BATCH_SUPPORT 121
#define SQL_CATALOG_LOCATION SQL_QUALIFIER_LOCATION
#define SQL_CATALOG_NAME_SEPARATOR SQL_QUALIFIER_NAME_SEPARATOR
#define SQL_CATALOG_TERM SQL_QUALIFIER_TERM
#define SQL_CATALOG_USAGE SQL_QUALIFIER_USAGE
#define SQL_CONVERT_WCHAR 122
#define SQL_CONVERT_INTERVAL_DAY_TIME 123
#define SQL_CONVERT_INTERVAL_YEAR_MONTH 124
#define SQL_CONVERT_WLONGVARCHAR 125
#define SQL_CONVERT_WVARCHAR 126
#define SQL_CREATE_ASSERTION 127
#define SQL_CREATE_CHARACTER_SET 128
#define SQL_CREATE_COLLATION 129
#define SQL_CREATE_DOMAIN 130
#define SQL_CREATE_SCHEMA 131
#define SQL_CREATE_TABLE 132
#define SQL_CREATE_TRANSLATION 133
#define SQL_CREATE_VIEW 134
#define SQL_DRIVER_HDESC 135
#define SQL_DROP_ASSERTION 136
#define SQL_DROP_CHARACTER_SET 137
#define SQL_DROP_COLLATION 138
#define SQL_DROP_DOMAIN 139
#define SQL_DROP_SCHEMA 140
#define SQL_DROP_TABLE 141
#define SQL_DROP_TRANSLATION 142
#define SQL_DROP_VIEW 143
#define SQL_DYNAMIC_CURSOR_ATTRIBUTES1 144
#define SQL_DYNAMIC_CURSOR_ATTRIBUTES2 145
#define SQL_FORWARD_ONLY_CURSOR_ATTRIBUTES1 146
#define SQL_FORWARD_ONLY_CURSOR_ATTRIBUTES2 147
#define SQL_INDEX_KEYWORDS 148
#define SQL_INFO_SCHEMA_VIEWS 149
#define SQL_KEYSET_CURSOR_ATTRIBUTES1 150
#define SQL_KEYSET_CURSOR_ATTRIBUTES2 151
#define SQL_MAX_ASYNC_CONCURRENT_STATEMENTS 10022 
#define SQL_ODBC_INTERFACE_CONFORMANCE 152
#define SQL_PARAM_ARRAY_ROW_COUNTS 153
#define SQL_PARAM_ARRAY_SELECTS 154
#define SQL_SCHEMA_TERM SQL_OWNER_TERM
#define SQL_SCHEMA_USAGE SQL_OWNER_USAGE
#define SQL_SQL92_DATETIME_FUNCTIONS 155
#define SQL_SQL92_FOREIGN_KEY_DELETE_RULE 156
#define SQL_SQL92_FOREIGN_KEY_UPDATE_RULE 157
#define SQL_SQL92_GRANT 158
#define SQL_SQL92_NUMERIC_VALUE_FUNCTIONS 159
#define SQL_SQL92_PREDICATES 160
#define SQL_SQL92_RELATIONAL_JOIN_OPERATORS 161
#define SQL_SQL92_REVOKE 162
#define SQL_SQL92_ROW_VALUE_CONSTRUCTOR 163
#define SQL_SQL92_STRING_FUNCTIONS 164
#define SQL_SQL92_VALUE_EXPRESSIONS 165
#define SQL_STANDARD_CLI_CONFORMANCE 166
#define SQL_STATIC_CURSOR_ATTRIBUTES1 167
#define SQL_STATIC_CURSOR_ATTRIBUTES2 168
#define SQL_AGGREGATE_FUNCTIONS 169
#define SQL_DDL_INDEX 170
#define SQL_DM_VER 171
#define SQL_INSERT_STATEMENT 172
#define SQL_CONVERT_GUID 173
#define SQL_UNION_STATEMENT SQL_UNION
#define SQL_DTC_TRANSITION_COST 1750
#define SQL_AT_ADD_COLUMN_SINGLE 0x00000020L
#define SQL_AT_ADD_COLUMN_DEFAULT 0x00000040L
#define SQL_AT_ADD_COLUMN_COLLATION 0x00000080L
#define SQL_AT_SET_COLUMN_DEFAULT 0x00000100L
#define SQL_AT_DROP_COLUMN_DEFAULT 0x00000200L
#define SQL_AT_DROP_COLUMN_CASCADE 0x00000400L
#define SQL_AT_DROP_COLUMN_RESTRICT 0x00000800L
#define SQL_AT_ADD_TABLE_CONSTRAINT 0x00001000L
#define SQL_AT_DROP_TABLE_CONSTRAINT_CASCADE 0x00002000L
#define SQL_AT_DROP_TABLE_CONSTRAINT_RESTRICT 0x00004000L
#define SQL_AT_CONSTRAINT_NAME_DEFINITION 0x00008000L
#define SQL_AT_CONSTRAINT_INITIALLY_DEFERRED 0x00010000L
#define SQL_AT_CONSTRAINT_INITIALLY_IMMEDIATE 0x00020000L
#define SQL_AT_CONSTRAINT_DEFERRABLE 0x00040000L
#define SQL_AT_CONSTRAINT_NON_DEFERRABLE 0x00080000L
#define SQL_CVT_CHAR 0x00000001L
#define SQL_CVT_NUMERIC 0x00000002L
#define SQL_CVT_DECIMAL 0x00000004L
#define SQL_CVT_INTEGER 0x00000008L
#define SQL_CVT_SMALLINT 0x00000010L
#define SQL_CVT_FLOAT 0x00000020L
#define SQL_CVT_REAL 0x00000040L
#define SQL_CVT_DOUBLE 0x00000080L
#define SQL_CVT_VARCHAR 0x00000100L
#define SQL_CVT_LONGVARCHAR 0x00000200L
#define SQL_CVT_BINARY 0x00000400L
#define SQL_CVT_VARBINARY 0x00000800L
#define SQL_CVT_BIT 0x00001000L
#define SQL_CVT_TINYINT 0x00002000L
#define SQL_CVT_BIGINT 0x00004000L
#define SQL_CVT_DATE 0x00008000L
#define SQL_CVT_TIME 0x00010000L
#define SQL_CVT_TIMESTAMP 0x00020000L
#define SQL_CVT_LONGVARBINARY 0x00040000L
#define SQL_CVT_INTERVAL_YEAR_MONTH 0x00080000L
#define SQL_CVT_INTERVAL_DAY_TIME 0x00100000L
#define SQL_CVT_WCHAR 0x00200000L
#define SQL_CVT_WLONGVARCHAR 0x00400000L
#define SQL_CVT_WVARCHAR 0x00800000L
#define SQL_CVT_GUID 0x01000000L
#define SQL_FN_CVT_CONVERT 0x00000001L
#define SQL_FN_CVT_CAST 0x00000002L
#define SQL_FN_STR_CONCAT 0x00000001L
#define SQL_FN_STR_INSERT 0x00000002L
#define SQL_FN_STR_LEFT 0x00000004L
#define SQL_FN_STR_LTRIM 0x00000008L
#define SQL_FN_STR_LENGTH 0x00000010L
#define SQL_FN_STR_LOCATE 0x00000020L
#define SQL_FN_STR_LCASE 0x00000040L
#define SQL_FN_STR_REPEAT 0x00000080L
#define SQL_FN_STR_REPLACE 0x00000100L
#define SQL_FN_STR_RIGHT 0x00000200L
#define SQL_FN_STR_RTRIM 0x00000400L
#define SQL_FN_STR_SUBSTRING 0x00000800L
#define SQL_FN_STR_UCASE 0x00001000L
#define SQL_FN_STR_ASCII 0x00002000L
#define SQL_FN_STR_CHAR 0x00004000L
#define SQL_FN_STR_DIFFERENCE 0x00008000L
#define SQL_FN_STR_LOCATE_2 0x00010000L
#define SQL_FN_STR_SOUNDEX 0x00020000L
#define SQL_FN_STR_SPACE 0x00040000L
#define SQL_FN_STR_BIT_LENGTH 0x00080000L
#define SQL_FN_STR_CHAR_LENGTH 0x00100000L
#define SQL_FN_STR_CHARACTER_LENGTH 0x00200000L
#define SQL_FN_STR_OCTET_LENGTH 0x00400000L
#define SQL_FN_STR_POSITION 0x00800000L
#define SQL_SSF_CONVERT 0x00000001L
#define SQL_SSF_LOWER 0x00000002L
#define SQL_SSF_UPPER 0x00000004L
#define SQL_SSF_SUBSTRING 0x00000008L
#define SQL_SSF_TRANSLATE 0x00000010L
#define SQL_SSF_TRIM_BOTH 0x00000020L
#define SQL_SSF_TRIM_LEADING 0x00000040L
#define SQL_SSF_TRIM_TRAILING 0x00000080L
#define SQL_FN_NUM_ABS 0x00000001L
#define SQL_FN_NUM_ACOS 0x00000002L
#define SQL_FN_NUM_ASIN 0x00000004L
#define SQL_FN_NUM_ATAN 0x00000008L
#define SQL_FN_NUM_ATAN2 0x00000010L
#define SQL_FN_NUM_CEILING 0x00000020L
#define SQL_FN_NUM_COS 0x00000040L
#define SQL_FN_NUM_COT 0x00000080L
#define SQL_FN_NUM_EXP 0x00000100L
#define SQL_FN_NUM_FLOOR 0x00000200L
#define SQL_FN_NUM_LOG 0x00000400L
#define SQL_FN_NUM_MOD 0x00000800L
#define SQL_FN_NUM_SIGN 0x00001000L
#define SQL_FN_NUM_SIN 0x00002000L
#define SQL_FN_NUM_SQRT 0x00004000L
#define SQL_FN_NUM_TAN 0x00008000L
#define SQL_FN_NUM_PI 0x00010000L
#define SQL_FN_NUM_RAND 0x00020000L
#define SQL_FN_NUM_DEGREES 0x00040000L
#define SQL_FN_NUM_LOG10 0x00080000L
#define SQL_FN_NUM_POWER 0x00100000L
#define SQL_FN_NUM_RADIANS 0x00200000L
#define SQL_FN_NUM_ROUND 0x00400000L
#define SQL_FN_NUM_TRUNCATE 0x00800000L
#define SQL_SNVF_BIT_LENGTH 0x00000001L
#define SQL_SNVF_CHAR_LENGTH 0x00000002L
#define SQL_SNVF_CHARACTER_LENGTH 0x00000004L
#define SQL_SNVF_EXTRACT 0x00000008L
#define SQL_SNVF_OCTET_LENGTH 0x00000010L
#define SQL_SNVF_POSITION 0x00000020L
#define SQL_FN_TD_NOW 0x00000001L
#define SQL_FN_TD_CURDATE 0x00000002L
#define SQL_FN_TD_DAYOFMONTH 0x00000004L
#define SQL_FN_TD_DAYOFWEEK 0x00000008L
#define SQL_FN_TD_DAYOFYEAR 0x00000010L
#define SQL_FN_TD_MONTH 0x00000020L
#define SQL_FN_TD_QUARTER 0x00000040L
#define SQL_FN_TD_WEEK 0x00000080L
#define SQL_FN_TD_YEAR 0x00000100L
#define SQL_FN_TD_CURTIME 0x00000200L
#define SQL_FN_TD_HOUR 0x00000400L
#define SQL_FN_TD_MINUTE 0x00000800L
#define SQL_FN_TD_SECOND 0x00001000L
#define SQL_FN_TD_TIMESTAMPADD 0x00002000L
#define SQL_FN_TD_TIMESTAMPDIFF 0x00004000L
#define SQL_FN_TD_DAYNAME 0x00008000L
#define SQL_FN_TD_MONTHNAME 0x00010000L
#define SQL_FN_TD_CURRENT_DATE 0x00020000L
#define SQL_FN_TD_CURRENT_TIME 0x00040000L
#define SQL_FN_TD_CURRENT_TIMESTAMP 0x00080000L
#define SQL_FN_TD_EXTRACT 0x00100000L
#define SQL_SDF_CURRENT_DATE 0x00000001L
#define SQL_SDF_CURRENT_TIME 0x00000002L
#define SQL_SDF_CURRENT_TIMESTAMP 0x00000004L
#define SQL_FN_SYS_USERNAME 0x00000001L
#define SQL_FN_SYS_DBNAME 0x00000002L
#define SQL_FN_SYS_IFNULL 0x00000004L
#define SQL_FN_TSI_FRAC_SECOND 0x00000001L
#define SQL_FN_TSI_SECOND 0x00000002L
#define SQL_FN_TSI_MINUTE 0x00000004L
#define SQL_FN_TSI_HOUR 0x00000008L
#define SQL_FN_TSI_DAY 0x00000010L
#define SQL_FN_TSI_WEEK 0x00000020L
#define SQL_FN_TSI_MONTH 0x00000040L
#define SQL_FN_TSI_QUARTER 0x00000080L
#define SQL_FN_TSI_YEAR 0x00000100L
#define SQL_CA1_NEXT 0x00000001L
#define SQL_CA1_ABSOLUTE 0x00000002L
#define SQL_CA1_RELATIVE 0x00000004L
#define SQL_CA1_BOOKMARK 0x00000008L
#define SQL_CA1_LOCK_NO_CHANGE 0x00000040L
#define SQL_CA1_LOCK_EXCLUSIVE 0x00000080L
#define SQL_CA1_LOCK_UNLOCK 0x00000100L
#define SQL_CA1_POS_POSITION 0x00000200L
#define SQL_CA1_POS_UPDATE 0x00000400L
#define SQL_CA1_POS_DELETE 0x00000800L
#define SQL_CA1_POS_REFRESH 0x00001000L
#define SQL_CA1_POSITIONED_UPDATE 0x00002000L
#define SQL_CA1_POSITIONED_DELETE 0x00004000L
#define SQL_CA1_SELECT_FOR_UPDATE 0x00008000L
#define SQL_CA1_BULK_ADD 0x00010000L
#define SQL_CA1_BULK_UPDATE_BY_BOOKMARK 0x00020000L
#define SQL_CA1_BULK_DELETE_BY_BOOKMARK 0x00040000L
#define SQL_CA1_BULK_FETCH_BY_BOOKMARK 0x00080000L
#define SQL_CA2_READ_ONLY_CONCURRENCY 0x00000001L
#define SQL_CA2_LOCK_CONCURRENCY 0x00000002L
#define SQL_CA2_OPT_ROWVER_CONCURRENCY 0x00000004L
#define SQL_CA2_OPT_VALUES_CONCURRENCY 0x00000008L
#define SQL_CA2_SENSITIVITY_ADDITIONS 0x00000010L
#define SQL_CA2_SENSITIVITY_DELETIONS 0x00000020L
#define SQL_CA2_SENSITIVITY_UPDATES 0x00000040L
#define SQL_CA2_MAX_ROWS_SELECT 0x00000080L
#define SQL_CA2_MAX_ROWS_INSERT 0x00000100L
#define SQL_CA2_MAX_ROWS_DELETE 0x00000200L
#define SQL_CA2_MAX_ROWS_UPDATE 0x00000400L
#define SQL_CA2_MAX_ROWS_CATALOG 0x00000800L
#define SQL_CA2_MAX_ROWS_AFFECTS_ALL 0xF80L
#define SQL_CA2_CRC_EXACT 0x00001000L
#define SQL_CA2_CRC_APPROXIMATE 0x00002000L
#define SQL_CA2_SIMULATE_NON_UNIQUE 0x00004000L
#define SQL_CA2_SIMULATE_TRY_UNIQUE 0x00008000L
#define SQL_CA2_SIMULATE_UNIQUE 0x00010000L
#define SQL_OAC_NONE 0x0000
#define SQL_OAC_LEVEL1 0x0001
#define SQL_OAC_LEVEL2 0x0002
#define SQL_OSCC_NOT_COMPLIANT 0x0000
#define SQL_OSCC_COMPLIANT 0x0001
#define SQL_OSC_MINIMUM 0x0000
#define SQL_OSC_CORE 0x0001
#define SQL_OSC_EXTENDED 0x0002
#define SQL_CB_NULL 0x0000
#define SQL_CB_NON_NULL 0x0001
#define SQL_SO_FORWARD_ONLY 0x00000001L
#define SQL_SO_KEYSET_DRIVEN 0x00000002L
#define SQL_SO_DYNAMIC 0x00000004L
#define SQL_SO_MIXED 0x00000008L
#define SQL_SO_STATIC 0x00000010L
#define SQL_FD_FETCH_RESUME 0x00000040L
#define SQL_FD_FETCH_BOOKMARK 0x00000080L
#define SQL_TXN_VERSIONING 0x00000010L
#define SQL_CN_NONE 0x0000
#define SQL_CN_DIFFERENT 0x0001
#define SQL_CN_ANY 0x0002
#define SQL_NNC_NULL 0x0000
#define SQL_NNC_NON_NULL 0x0001
#define SQL_NC_START 0x0002
#define SQL_NC_END 0x0004
#define SQL_FILE_NOT_SUPPORTED 0x0000
#define SQL_FILE_TABLE 0x0001
#define SQL_FILE_QUALIFIER 0x0002
#define SQL_FILE_CATALOG SQL_FILE_QUALIFIER
#define SQL_GD_BLOCK 0x00000004L
#define SQL_GD_BOUND 0x00000008L
#define SQL_PS_POSITIONED_DELETE 0x00000001L
#define SQL_PS_POSITIONED_UPDATE 0x00000002L
#define SQL_PS_SELECT_FOR_UPDATE 0x00000004L
#define SQL_GB_NOT_SUPPORTED 0x0000
#define SQL_GB_GROUP_BY_EQUALS_SELECT 0x0001
#define SQL_GB_GROUP_BY_CONTAINS_SELECT 0x0002
#define SQL_GB_NO_RELATION 0x0003
#define SQL_GB_COLLATE 0x0004
#define SQL_OU_DML_STATEMENTS 0x00000001L
#define SQL_OU_PROCEDURE_INVOCATION 0x00000002L
#define SQL_OU_TABLE_DEFINITION 0x00000004L
#define SQL_OU_INDEX_DEFINITION 0x00000008L
#define SQL_OU_PRIVILEGE_DEFINITION 0x00000010L
#define SQL_SU_DML_STATEMENTS SQL_OU_DML_STATEMENTS
#define SQL_SU_PROCEDURE_INVOCATION SQL_OU_PROCEDURE_INVOCATION
#define SQL_SU_TABLE_DEFINITION SQL_OU_TABLE_DEFINITION
#define SQL_SU_INDEX_DEFINITION SQL_OU_INDEX_DEFINITION
#define SQL_SU_PRIVILEGE_DEFINITION SQL_OU_PRIVILEGE_DEFINITION
#define SQL_QU_DML_STATEMENTS 0x00000001L
#define SQL_QU_PROCEDURE_INVOCATION 0x00000002L
#define SQL_QU_TABLE_DEFINITION 0x00000004L
#define SQL_QU_INDEX_DEFINITION 0x00000008L
#define SQL_QU_PRIVILEGE_DEFINITION 0x00000010L
#define SQL_CU_DML_STATEMENTS SQL_QU_DML_STATEMENTS
#define SQL_CU_PROCEDURE_INVOCATION SQL_QU_PROCEDURE_INVOCATION
#define SQL_CU_TABLE_DEFINITION SQL_QU_TABLE_DEFINITION
#define SQL_CU_INDEX_DEFINITION SQL_QU_INDEX_DEFINITION
#define SQL_CU_PRIVILEGE_DEFINITION SQL_QU_PRIVILEGE_DEFINITION
#define SQL_SQ_COMPARISON 0x00000001L
#define SQL_SQ_EXISTS 0x00000002L
#define SQL_SQ_IN 0x00000004L
#define SQL_SQ_QUANTIFIED 0x00000008L
#define SQL_SQ_CORRELATED_SUBQUERIES 0x00000010L
#define SQL_U_UNION 0x00000001L
#define SQL_U_UNION_ALL 0x00000002L
#define SQL_BP_CLOSE 0x00000001L
#define SQL_BP_DELETE 0x00000002L
#define SQL_BP_DROP 0x00000004L
#define SQL_BP_TRANSACTION 0x00000008L
#define SQL_BP_UPDATE 0x00000010L
#define SQL_BP_OTHER_HSTMT 0x00000020L
#define SQL_BP_SCROLL 0x00000040L
#define SQL_SS_ADDITIONS 0x00000001L
#define SQL_SS_DELETIONS 0x00000002L
#define SQL_SS_UPDATES 0x00000004L
#define SQL_CV_CREATE_VIEW 0x00000001L
#define SQL_CV_CHECK_OPTION 0x00000002L
#define SQL_CV_CASCADED 0x00000004L
#define SQL_CV_LOCAL 0x00000008L
#define SQL_LCK_NO_CHANGE 0x00000001L
#define SQL_LCK_EXCLUSIVE 0x00000002L
#define SQL_LCK_UNLOCK 0x00000004L
#define SQL_POS_POSITION 0x00000001L
#define SQL_POS_REFRESH 0x00000002L
#define SQL_POS_UPDATE 0x00000004L
#define SQL_POS_DELETE 0x00000008L
#define SQL_POS_ADD 0x00000010L
#define SQL_QL_START 0x0001
#define SQL_QL_END 0x0002
#define SQL_AF_AVG 0x00000001L
#define SQL_AF_COUNT 0x00000002L
#define SQL_AF_MAX 0x00000004L
#define SQL_AF_MIN 0x00000008L
#define SQL_AF_SUM 0x00000010L
#define SQL_AF_DISTINCT 0x00000020L
#define SQL_AF_ALL 0x00000040L
#define SQL_SC_SQL92_ENTRY 0x00000001L
#define SQL_SC_FIPS127_2_TRANSITIONAL 0x00000002L
#define SQL_SC_SQL92_INTERMEDIATE 0x00000004L
#define SQL_SC_SQL92_FULL 0x00000008L
#define SQL_DL_SQL92_DATE 0x00000001L
#define SQL_DL_SQL92_TIME 0x00000002L
#define SQL_DL_SQL92_TIMESTAMP 0x00000004L
#define SQL_DL_SQL92_INTERVAL_YEAR 0x00000008L
#define SQL_DL_SQL92_INTERVAL_MONTH 0x00000010L
#define SQL_DL_SQL92_INTERVAL_DAY 0x00000020L
#define SQL_DL_SQL92_INTERVAL_HOUR 0x00000040L
#define SQL_DL_SQL92_INTERVAL_MINUTE 0x00000080L
#define SQL_DL_SQL92_INTERVAL_SECOND 0x00000100L
#define SQL_DL_SQL92_INTERVAL_YEAR_TO_MONTH 0x00000200L
#define SQL_DL_SQL92_INTERVAL_DAY_TO_HOUR 0x00000400L
#define SQL_DL_SQL92_INTERVAL_DAY_TO_MINUTE 0x00000800L
#define SQL_DL_SQL92_INTERVAL_DAY_TO_SECOND 0x00001000L
#define SQL_DL_SQL92_INTERVAL_HOUR_TO_MINUTE 0x00002000L
#define SQL_DL_SQL92_INTERVAL_HOUR_TO_SECOND 0x00004000L
#define SQL_DL_SQL92_INTERVAL_MINUTE_TO_SECOND 0x00008000L
#define SQL_CL_START SQL_QL_START
#define SQL_CL_END SQL_QL_END
#define SQL_BRC_PROCEDURES 0x0000001
#define SQL_BRC_EXPLICIT 0x0000002
#define SQL_BRC_ROLLED_UP 0x0000004
#define SQL_BS_SELECT_EXPLICIT 0x00000001L
#define SQL_BS_ROW_COUNT_EXPLICIT 0x00000002L
#define SQL_BS_SELECT_PROC 0x00000004L
#define SQL_BS_ROW_COUNT_PROC 0x00000008L
#define SQL_PARC_BATCH 1
#define SQL_PARC_NO_BATCH 2
#define SQL_PAS_BATCH 1
#define SQL_PAS_NO_BATCH 2
#define SQL_PAS_NO_SELECT 3
#define SQL_IK_NONE 0x00000000L
#define SQL_IK_ASC 0x00000001L
#define SQL_IK_DESC 0x00000002L
#define SQL_IK_ALL 0x00000003L
#define SQL_ISV_ASSERTIONS 0x00000001L
#define SQL_ISV_CHARACTER_SETS 0x00000002L
#define SQL_ISV_CHECK_CONSTRAINTS 0x00000004L
#define SQL_ISV_COLLATIONS 0x00000008L
#define SQL_ISV_COLUMN_DOMAIN_USAGE 0x00000010L
#define SQL_ISV_COLUMN_PRIVILEGES 0x00000020L
#define SQL_ISV_COLUMNS 0x00000040L
#define SQL_ISV_CONSTRAINT_COLUMN_USAGE 0x00000080L
#define SQL_ISV_CONSTRAINT_TABLE_USAGE 0x00000100L
#define SQL_ISV_DOMAIN_CONSTRAINTS 0x00000200L
#define SQL_ISV_DOMAINS 0x00000400L
#define SQL_ISV_KEY_COLUMN_USAGE 0x00000800L
#define SQL_ISV_REFERENTIAL_CONSTRAINTS 0x00001000L
#define SQL_ISV_SCHEMATA 0x00002000L
#define SQL_ISV_SQL_LANGUAGES 0x00004000L
#define SQL_ISV_TABLE_CONSTRAINTS 0x00008000L
#define SQL_ISV_TABLE_PRIVILEGES 0x00010000L
#define SQL_ISV_TABLES 0x00020000L
#define SQL_ISV_TRANSLATIONS 0x00040000L
#define SQL_ISV_USAGE_PRIVILEGES 0x00080000L
#define SQL_ISV_VIEW_COLUMN_USAGE 0x00100000L
#define SQL_ISV_VIEW_TABLE_USAGE 0x00200000L
#define SQL_ISV_VIEWS 0x00400000L
#define SQL_AD_CONSTRAINT_NAME_DEFINITION 0x00000001L
#define SQL_AD_ADD_DOMAIN_CONSTRAINT 0x00000002L
#define SQL_AD_DROP_DOMAIN_CONSTRAINT 0x00000004L
#define SQL_AD_ADD_DOMAIN_DEFAULT 0x00000008L
#define SQL_AD_DROP_DOMAIN_DEFAULT 0x00000010L
#define SQL_AD_ADD_CONSTRAINT_INITIALLY_DEFERRED 0x00000020L
#define SQL_AD_ADD_CONSTRAINT_INITIALLY_IMMEDIATE 0x00000040L
#define SQL_AD_ADD_CONSTRAINT_DEFERRABLE 0x00000080L
#define SQL_AD_ADD_CONSTRAINT_NON_DEFERRABLE 0x00000100L
#define SQL_CS_CREATE_SCHEMA 0x00000001L
#define SQL_CS_AUTHORIZATION 0x00000002L
#define SQL_CS_DEFAULT_CHARACTER_SET 0x00000004L
#define SQL_CTR_CREATE_TRANSLATION 0x00000001L
#define SQL_CA_CREATE_ASSERTION 0x00000001L
#define SQL_CA_CONSTRAINT_INITIALLY_DEFERRED 0x00000010L
#define SQL_CA_CONSTRAINT_INITIALLY_IMMEDIATE 0x00000020L
#define SQL_CA_CONSTRAINT_DEFERRABLE 0x00000040L
#define SQL_CA_CONSTRAINT_NON_DEFERRABLE 0x00000080L
#define SQL_CCS_CREATE_CHARACTER_SET 0x00000001L
#define SQL_CCS_COLLATE_CLAUSE 0x00000002L
#define SQL_CCS_LIMITED_COLLATION 0x00000004L
#define SQL_CCOL_CREATE_COLLATION 0x00000001L
#define SQL_CDO_CREATE_DOMAIN 0x00000001L
#define SQL_CDO_DEFAULT 0x00000002L
#define SQL_CDO_CONSTRAINT 0x00000004L
#define SQL_CDO_COLLATION 0x00000008L
#define SQL_CDO_CONSTRAINT_NAME_DEFINITION 0x00000010L
#define SQL_CDO_CONSTRAINT_INITIALLY_DEFERRED 0x00000020L
#define SQL_CDO_CONSTRAINT_INITIALLY_IMMEDIATE 0x00000040L
#define SQL_CDO_CONSTRAINT_DEFERRABLE 0x00000080L
#define SQL_CDO_CONSTRAINT_NON_DEFERRABLE 0x00000100L
#define SQL_CT_CREATE_TABLE 0x00000001L
#define SQL_CT_COMMIT_PRESERVE 0x00000002L
#define SQL_CT_COMMIT_DELETE 0x00000004L
#define SQL_CT_GLOBAL_TEMPORARY 0x00000008L
#define SQL_CT_LOCAL_TEMPORARY 0x00000010L
#define SQL_CT_CONSTRAINT_INITIALLY_DEFERRED 0x00000020L
#define SQL_CT_CONSTRAINT_INITIALLY_IMMEDIATE 0x00000040L
#define SQL_CT_CONSTRAINT_DEFERRABLE 0x00000080L
#define SQL_CT_CONSTRAINT_NON_DEFERRABLE 0x00000100L
#define SQL_CT_COLUMN_CONSTRAINT 0x00000200L
#define SQL_CT_COLUMN_DEFAULT 0x00000400L
#define SQL_CT_COLUMN_COLLATION 0x00000800L
#define SQL_CT_TABLE_CONSTRAINT 0x00001000L
#define SQL_CT_CONSTRAINT_NAME_DEFINITION 0x00002000L
#define SQL_DI_CREATE_INDEX 0x00000001L
#define SQL_DI_DROP_INDEX 0x00000002L
#define SQL_DC_DROP_COLLATION 0x00000001L
#define SQL_DD_DROP_DOMAIN 0x00000001L
#define SQL_DD_RESTRICT 0x00000002L
#define SQL_DD_CASCADE 0x00000004L
#define SQL_DS_DROP_SCHEMA 0x00000001L
#define SQL_DS_RESTRICT 0x00000002L
#define SQL_DS_CASCADE 0x00000004L
#define SQL_DCS_DROP_CHARACTER_SET 0x00000001L
#define SQL_DA_DROP_ASSERTION 0x00000001L
#define SQL_DT_DROP_TABLE 0x00000001L
#define SQL_DT_RESTRICT 0x00000002L
#define SQL_DT_CASCADE 0x00000004L
#define SQL_DTR_DROP_TRANSLATION 0x00000001L
#define SQL_DV_DROP_VIEW 0x00000001L
#define SQL_DV_RESTRICT 0x00000002L
#define SQL_DV_CASCADE 0x00000004L
#define SQL_IS_INSERT_LITERALS 0x00000001L
#define SQL_IS_INSERT_SEARCHED 0x00000002L
#define SQL_IS_SELECT_INTO 0x00000004L
#define SQL_OIC_CORE 1U
#define SQL_OIC_LEVEL1 2U
#define SQL_OIC_LEVEL2 3U
#define SQL_SFKD_CASCADE 0x00000001L
#define SQL_SFKD_NO_ACTION 0x00000002L
#define SQL_SFKD_SET_DEFAULT 0x00000004L
#define SQL_SFKD_SET_NULL 0x00000008L
#define SQL_SFKU_CASCADE 0x00000001L
#define SQL_SFKU_NO_ACTION 0x00000002L
#define SQL_SFKU_SET_DEFAULT 0x00000004L
#define SQL_SFKU_SET_NULL 0x00000008L
#define SQL_SG_USAGE_ON_DOMAIN 0x00000001L
#define SQL_SG_USAGE_ON_CHARACTER_SET 0x00000002L
#define SQL_SG_USAGE_ON_COLLATION 0x00000004L
#define SQL_SG_USAGE_ON_TRANSLATION 0x00000008L
#define SQL_SG_WITH_GRANT_OPTION 0x00000010L
#define SQL_SG_DELETE_TABLE 0x00000020L
#define SQL_SG_INSERT_TABLE 0x00000040L
#define SQL_SG_INSERT_COLUMN 0x00000080L
#define SQL_SG_REFERENCES_TABLE 0x00000100L
#define SQL_SG_REFERENCES_COLUMN 0x00000200L
#define SQL_SG_SELECT_TABLE 0x00000400L
#define SQL_SG_UPDATE_TABLE 0x00000800L
#define SQL_SG_UPDATE_COLUMN 0x00001000L
#define SQL_SP_EXISTS 0x00000001L
#define SQL_SP_ISNOTNULL 0x00000002L
#define SQL_SP_ISNULL 0x00000004L
#define SQL_SP_MATCH_FULL 0x00000008L
#define SQL_SP_MATCH_PARTIAL 0x00000010L
#define SQL_SP_MATCH_UNIQUE_FULL 0x00000020L
#define SQL_SP_MATCH_UNIQUE_PARTIAL 0x00000040L
#define SQL_SP_OVERLAPS 0x00000080L
#define SQL_SP_UNIQUE 0x00000100L
#define SQL_SP_LIKE 0x00000200L
#define SQL_SP_IN 0x00000400L
#define SQL_SP_BETWEEN 0x00000800L
#define SQL_SP_COMPARISON 0x00001000L
#define SQL_SP_QUANTIFIED_COMPARISON 0x00002000L
#define SQL_SRJO_CORRESPONDING_CLAUSE 0x00000001L
#define SQL_SRJO_CROSS_JOIN 0x00000002L
#define SQL_SRJO_EXCEPT_JOIN 0x00000004L
#define SQL_SRJO_FULL_OUTER_JOIN 0x00000008L
#define SQL_SRJO_INNER_JOIN 0x00000010L
#define SQL_SRJO_INTERSECT_JOIN 0x00000020L
#define SQL_SRJO_LEFT_OUTER_JOIN 0x00000040L
#define SQL_SRJO_NATURAL_JOIN 0x00000080L
#define SQL_SRJO_RIGHT_OUTER_JOIN 0x00000100L
#define SQL_SRJO_UNION_JOIN 0x00000200L
#define SQL_SR_USAGE_ON_DOMAIN 0x00000001L
#define SQL_SR_USAGE_ON_CHARACTER_SET 0x00000002L
#define SQL_SR_USAGE_ON_COLLATION 0x00000004L
#define SQL_SR_USAGE_ON_TRANSLATION 0x00000008L
#define SQL_SR_GRANT_OPTION_FOR 0x00000010L
#define SQL_SR_CASCADE 0x00000020L
#define SQL_SR_RESTRICT 0x00000040L
#define SQL_SR_DELETE_TABLE 0x00000080L
#define SQL_SR_INSERT_TABLE 0x00000100L
#define SQL_SR_INSERT_COLUMN 0x00000200L
#define SQL_SR_REFERENCES_TABLE 0x00000400L
#define SQL_SR_REFERENCES_COLUMN 0x00000800L
#define SQL_SR_SELECT_TABLE 0x00001000L
#define SQL_SR_UPDATE_TABLE 0x00002000L
#define SQL_SR_UPDATE_COLUMN 0x00004000L
#define SQL_SRVC_VALUE_EXPRESSION 0x00000001L
#define SQL_SRVC_NULL 0x00000002L
#define SQL_SRVC_DEFAULT 0x00000004L
#define SQL_SRVC_ROW_SUBQUERY 0x00000008L
#define SQL_SVE_CASE 0x00000001L
#define SQL_SVE_CAST 0x00000002L
#define SQL_SVE_COALESCE 0x00000004L
#define SQL_SVE_NULLIF 0x00000008L
#define SQL_SCC_XOPEN_CLI_VERSION1 0x00000001L
#define SQL_SCC_ISO92_CLI 0x00000002L
#define SQL_US_UNION SQL_U_UNION
#define SQL_US_UNION_ALL SQL_U_UNION_ALL
#define SQL_DTC_ENLIST_EXPENSIVE 0x00000001L
#define SQL_DTC_UNENLIST_EXPENSIVE 0x00000002L
#define SQL_FETCH_FIRST_USER 31
#define SQL_FETCH_FIRST_SYSTEM 32
#define SQL_ENTIRE_ROWSET 0
#define SQL_POSITION 0 
#define SQL_REFRESH 1 
#define SQL_UPDATE 2
#define SQL_DELETE 3
#define SQL_ADD 4
#define SQL_SETPOS_MAX_OPTION_VALUE SQL_ADD
#define SQL_UPDATE_BY_BOOKMARK 5
#define SQL_DELETE_BY_BOOKMARK 6
#define SQL_FETCH_BY_BOOKMARK 7
#define SQL_LOCK_NO_CHANGE 0 
#define SQL_LOCK_EXCLUSIVE 1 
#define SQL_LOCK_UNLOCK 2
#define SQL_SETPOS_MAX_LOCK_VALUE SQL_LOCK_UNLOCK
#define SQL_BEST_ROWID 1
#define SQL_ROWVER 2
#define SQL_PC_NOT_PSEUDO 1
#define SQL_QUICK 0
#define SQL_ENSURE 1
#define SQL_TABLE_STAT 0
#define SQL_ALL_CATALOGS "%"
#define SQL_ALL_SCHEMAS "%"
#define SQL_ALL_TABLE_TYPES "%"
#define SQL_DRIVER_NOPROMPT 0
#define SQL_DRIVER_COMPLETE 1
#define SQL_DRIVER_PROMPT 2
#define SQL_DRIVER_COMPLETE_REQUIRED 3
#define SQL_FETCH_BOOKMARK 8
#define SQL_ROW_SUCCESS 0
#define SQL_ROW_DELETED 1
#define SQL_ROW_UPDATED 2
#define SQL_ROW_NOROW 3
#define SQL_ROW_ADDED 4
#define SQL_ROW_ERROR 5
#define SQL_ROW_SUCCESS_WITH_INFO 6
#define SQL_ROW_PROCEED 0
#define SQL_ROW_IGNORE 1
#define SQL_PARAM_SUCCESS 0
#define SQL_PARAM_SUCCESS_WITH_INFO 6
#define SQL_PARAM_ERROR 5
#define SQL_PARAM_UNUSED 7
#define SQL_PARAM_DIAG_UNAVAILABLE 1
#define SQL_PARAM_PROCEED 0
#define SQL_PARAM_IGNORE 1
#define SQL_CASCADE 0
#define SQL_RESTRICT 1
#define SQL_SET_NULL 2
#define SQL_NO_ACTION 3
#define SQL_SET_DEFAULT 4
#define SQL_INITIALLY_DEFERRED 5
#define SQL_INITIALLY_IMMEDIATE 6
#define SQL_NOT_DEFERRABLE 7
#define SQL_PARAM_TYPE_UNKNOWN 0
#define SQL_PARAM_INPUT 1
#define SQL_RESULT_COL 3
#define SQL_PARAM_OUTPUT 4
#define SQL_RETURN_VALUE 5
#define SQL_PT_UNKNOWN 0
#define SQL_PT_PROCEDURE 1
#define SQL_PT_FUNCTION 2
#define SQL_DATABASE_NAME 16 
#define SQL_FD_FETCH_PREV SQL_FD_FETCH_PRIOR
#define SQL_FETCH_PREV SQL_FETCH_PRIOR
#define SQL_CONCUR_TIMESTAMP SQL_CONCUR_ROWVER
#define SQL_SCCO_OPT_TIMESTAMP SQL_SCCO_OPT_ROWVER
#define SQL_CC_DELETE SQL_CB_DELETE
#define SQL_CR_DELETE SQL_CB_DELETE
#define SQL_CC_CLOSE SQL_CB_CLOSE
#define SQL_CR_CLOSE SQL_CB_CLOSE
#define SQL_CC_PRESERVE SQL_CB_PRESERVE
#define SQL_CR_PRESERVE SQL_CB_PRESERVE
#define SQL_FETCH_RESUME 7
#define SQL_SCROLL_FORWARD_ONLY 0L 
#define SQL_SCROLL_KEYSET_DRIVEN (-1L) 
#define SQL_SCROLL_DYNAMIC (-2L) 
#define SQL_SCROLL_STATIC (-3L) 
#define TRACE_VERSION 1000 
#define TRACE_ON 0x00000001L
#define TRACE_VS_EVENT_ON 0x00000002L
#define ODBC_VS_FLAG_UNICODE_ARG 0x00000001L 
#define ODBC_VS_FLAG_UNICODE_COR 0x00000002L 
#define ODBC_VS_FLAG_RETCODE 0x00000004L 
#define ODBC_VS_FLAG_STOP 0x00000008L 
#define SQL_C_WCHAR SQL_WCHAR
#define SQL_C_TCHAR SQL_C_CHAR
#define SQL_SQLSTATE_SIZEW 10 
#define LINE_ADDRESSSTATE 0L
#define LINE_CALLINFO 1L
#define LINE_CALLSTATE 2L
#define LINE_CLOSE 3L
#define LINE_DEVSPECIFIC 4L
#define LINE_DEVSPECIFICFEATURE 5L
#define LINE_GATHERDIGITS 6L
#define LINE_GENERATE 7L
#define LINE_LINEDEVSTATE 8L
#define LINE_MONITORDIGITS 9L
#define LINE_MONITORMEDIA 10L
#define LINE_MONITORTONE 11L
#define LINE_REPLY 12L
#define LINE_REQUEST 13L
#define PHONE_BUTTON 14L
#define PHONE_CLOSE 15L
#define PHONE_DEVSPECIFIC 16L
#define PHONE_REPLY 17L
#define PHONE_STATE 18L
#define LINE_CREATE 19L
#define PHONE_CREATE 20L
#define TAPI_REPLY WM_USER + 99
#define TAPIERR_CONNECTED 0L
#define TAPIERR_DROPPED -1L
#define TAPIERR_NOREQUESTRECIPIENT -2L
#define TAPIERR_REQUESTQUEUEFULL -3L
#define TAPIERR_INVALDESTADDRESS -4L
#define TAPIERR_INVALWINDOWHANDLE -5L
#define TAPIERR_INVALDEVICECLASS -6L
#define TAPIERR_INVALDEVICEID -7L
#define TAPIERR_DEVICECLASSUNAVAIL -8L
#define TAPIERR_DEVICEIDUNAVAIL -9L
#define TAPIERR_DEVICEINUSE -10L
#define TAPIERR_DESTBUSY -11L
#define TAPIERR_DESTNOANSWER -12L
#define TAPIERR_DESTUNAVAIL -13L
#define TAPIERR_UNKNOWNWINHANDLE -14L
#define TAPIERR_UNKNOWNREQUESTID -15L
#define TAPIERR_REQUESTFAILED -16L
#define TAPIERR_REQUESTCANCELLED -17L
#define TAPIERR_INVALPOINTER -18L
#define TAPIMAXDESTADDRESSSIZE 80L
#define TAPIMAXAPPNAMESIZE 40L
#define TAPIMAXCALLEDPARTYSIZE 40L
#define TAPIMAXCOMMENTSIZE 80L
#define TAPIMAXDEVICECLASSSIZE 40L
#define TAPIMAXDEVICEIDSIZE 40L
#define PHONEBUTTONFUNCTION_UNKNOWN 0x00000000
#define PHONEBUTTONFUNCTION_CONFERENCE 0x00000001
#define PHONEBUTTONFUNCTION_TRANSFER 0x00000002
#define PHONEBUTTONFUNCTION_DROP 0x00000003
#define PHONEBUTTONFUNCTION_HOLD 0x00000004
#define PHONEBUTTONFUNCTION_RECALL 0x00000005
#define PHONEBUTTONFUNCTION_DISCONNECT 0x00000006
#define PHONEBUTTONFUNCTION_CONNECT 0x00000007
#define PHONEBUTTONFUNCTION_MSGWAITON 0x00000008
#define PHONEBUTTONFUNCTION_MSGWAITOFF 0x00000009
#define PHONEBUTTONFUNCTION_SELECTRING 0x0000000A
#define PHONEBUTTONFUNCTION_ABBREVDIAL 0x0000000B
#define PHONEBUTTONFUNCTION_FORWARD 0x0000000C
#define PHONEBUTTONFUNCTION_PICKUP 0x0000000D
#define PHONEBUTTONFUNCTION_RINGAGAIN 0x0000000E
#define PHONEBUTTONFUNCTION_PARK 0x0000000F
#define PHONEBUTTONFUNCTION_REJECT 0x00000010
#define PHONEBUTTONFUNCTION_REDIRECT 0x00000011
#define PHONEBUTTONFUNCTION_MUTE 0x00000012
#define PHONEBUTTONFUNCTION_VOLUMEUP 0x00000013
#define PHONEBUTTONFUNCTION_VOLUMEDOWN 0x00000014
#define PHONEBUTTONFUNCTION_SPEAKERON 0x00000015
#define PHONEBUTTONFUNCTION_SPEAKEROFF 0x00000016
#define PHONEBUTTONFUNCTION_FLASH 0x00000017
#define PHONEBUTTONFUNCTION_DATAON 0x00000018
#define PHONEBUTTONFUNCTION_DATAOFF 0x00000019
#define PHONEBUTTONFUNCTION_DONOTDISTURB 0x0000001A
#define PHONEBUTTONFUNCTION_INTERCOM 0x0000001B
#define PHONEBUTTONFUNCTION_BRIDGEDAPP 0x0000001C
#define PHONEBUTTONFUNCTION_BUSY 0x0000001D
#define PHONEBUTTONFUNCTION_CALLAPP 0x0000001E
#define PHONEBUTTONFUNCTION_DATETIME 0x0000001F
#define PHONEBUTTONFUNCTION_DIRECTORY 0x00000020
#define PHONEBUTTONFUNCTION_COVER 0x00000021
#define PHONEBUTTONFUNCTION_CALLID 0x00000022
#define PHONEBUTTONFUNCTION_LASTNUM 0x00000023
#define PHONEBUTTONFUNCTION_NIGHTSRV 0x00000024
#define PHONEBUTTONFUNCTION_SENDCALLS 0x00000025
#define PHONEBUTTONFUNCTION_MSGINDICATOR 0x00000026
#define PHONEBUTTONFUNCTION_REPDIAL 0x00000027
#define PHONEBUTTONFUNCTION_SETREPDIAL 0x00000028
#define PHONEBUTTONFUNCTION_SYSTEMSPEED 0x00000029
#define PHONEBUTTONFUNCTION_STATIONSPEED 0x0000002A
#define PHONEBUTTONFUNCTION_CAMPON 0x0000002B
#define PHONEBUTTONFUNCTION_SAVEREPEAT 0x0000002C
#define PHONEBUTTONFUNCTION_QUEUECALL 0x0000002D
#define PHONEBUTTONFUNCTION_NONE 0x0000002E
#define PHONEBUTTONMODE_DUMMY 0x00000001
#define PHONEBUTTONMODE_CALL 0x00000002
#define PHONEBUTTONMODE_FEATURE 0x00000004
#define PHONEBUTTONMODE_KEYPAD 0x00000008
#define PHONEBUTTONMODE_LOCAL 0x00000010
#define PHONEBUTTONMODE_DISPLAY 0x00000020
#define PHONEBUTTONSTATE_UP 0x00000001
#define PHONEBUTTONSTATE_DOWN 0x00000002
#define PHONEBUTTONSTATE_UNKNOWN 0x00000004
#define PHONEBUTTONSTATE_UNAVAIL 0x00000008
#define PHONEERR_ALLOCATED 0x90000001
#define PHONEERR_BADDEVICEID 0x90000002
#define PHONEERR_INCOMPATIBLEAPIVERSION 0x90000003
#define PHONEERR_INCOMPATIBLEEXTVERSION 0x90000004
#define PHONEERR_INIFILECORRUPT 0x90000005
#define PHONEERR_INUSE 0x90000006
#define PHONEERR_INVALAPPHANDLE 0x90000007
#define PHONEERR_INVALAPPNAME 0x90000008
#define PHONEERR_INVALBUTTONLAMPID 0x90000009
#define PHONEERR_INVALBUTTONMODE 0x9000000A
#define PHONEERR_INVALBUTTONSTATE 0x9000000B
#define PHONEERR_INVALDATAID 0x9000000C
#define PHONEERR_INVALDEVICECLASS 0x9000000D
#define PHONEERR_INVALEXTVERSION 0x9000000E
#define PHONEERR_INVALHOOKSWITCHDEV 0x9000000F
#define PHONEERR_INVALHOOKSWITCHMODE 0x90000010
#define PHONEERR_INVALLAMPMODE 0x90000011
#define PHONEERR_INVALPARAM 0x90000012
#define PHONEERR_INVALPHONEHANDLE 0x90000013
#define PHONEERR_INVALPHONESTATE 0x90000014
#define PHONEERR_INVALPOINTER 0x90000015
#define PHONEERR_INVALPRIVILEGE 0x90000016
#define PHONEERR_INVALRINGMODE 0x90000017
#define PHONEERR_NODEVICE 0x90000018
#define PHONEERR_NODRIVER 0x90000019
#define PHONEERR_NOMEM 0x9000001A
#define PHONEERR_NOTOWNER 0x9000001B
#define PHONEERR_OPERATIONFAILED 0x9000001C
#define PHONEERR_OPERATIONUNAVAIL 0x9000001D
#define PHONEERR_RESOURCEUNAVAIL 0x9000001F
#define PHONEERR_REQUESTOVERRUN 0x90000020
#define PHONEERR_STRUCTURETOOSMALL 0x90000021
#define PHONEERR_UNINITIALIZED 0x90000022
#define PHONEERR_REINIT 0x90000023
#define PHONEHOOKSWITCHDEV_HANDSET 0x00000001
#define PHONEHOOKSWITCHDEV_SPEAKER 0x00000002
#define PHONEHOOKSWITCHDEV_HEADSET 0x00000004
#define PHONEHOOKSWITCHMODE_ONHOOK 0x00000001
#define PHONEHOOKSWITCHMODE_MIC 0x00000002
#define PHONEHOOKSWITCHMODE_SPEAKER 0x00000004
#define PHONEHOOKSWITCHMODE_MICSPEAKER 0x00000008
#define PHONEHOOKSWITCHMODE_UNKNOWN 0x00000010
#define PHONELAMPMODE_DUMMY 0x00000001
#define PHONELAMPMODE_OFF 0x00000002
#define PHONELAMPMODE_STEADY 0x00000004
#define PHONELAMPMODE_WINK 0x00000008
#define PHONELAMPMODE_FLASH 0x00000010
#define PHONELAMPMODE_FLUTTER 0x00000020
#define PHONELAMPMODE_BROKENFLUTTER 0x00000040
#define PHONELAMPMODE_UNKNOWN 0x00000080
#define PHONEPRIVILEGE_MONITOR 0x00000001
#define PHONEPRIVILEGE_OWNER 0x00000002
#define PHONESTATE_OTHER 0x00000001
#define PHONESTATE_CONNECTED 0x00000002
#define PHONESTATE_DISCONNECTED 0x00000004
#define PHONESTATE_OWNER 0x00000008
#define PHONESTATE_MONITORS 0x00000010
#define PHONESTATE_DISPLAY 0x00000020
#define PHONESTATE_LAMP 0x00000040
#define PHONESTATE_RINGMODE 0x00000080
#define PHONESTATE_RINGVOLUME 0x00000100
#define PHONESTATE_HANDSETHOOKSWITCH 0x00000200
#define PHONESTATE_HANDSETVOLUME 0x00000400
#define PHONESTATE_HANDSETGAIN 0x00000800
#define PHONESTATE_SPEAKERHOOKSWITCH 0x00001000
#define PHONESTATE_SPEAKERVOLUME 0x00002000
#define PHONESTATE_SPEAKERGAIN 0x00004000
#define PHONESTATE_HEADSETHOOKSWITCH 0x00008000
#define PHONESTATE_HEADSETVOLUME 0x00010000
#define PHONESTATE_HEADSETGAIN 0x00020000
#define PHONESTATE_SUSPEND 0x00040000
#define PHONESTATE_RESUME 0x00080000
#define PHONESTATE_DEVSPECIFIC 0x00100000
#define PHONESTATE_REINIT 0x00200000
#define PHONESTATE_CAPSCHANGE 0x00400000
#define PHONESTATE_REMOVED 0x00800000
#define PHONESTATUSFLAGS_CONNECTED 0x00000001
#define PHONESTATUSFLAGS_SUSPENDED 0x00000002
#define STRINGFORMAT_ASCII 0x00000001
#define STRINGFORMAT_DBCS 0x00000002
#define STRINGFORMAT_UNICODE 0x00000003
#define STRINGFORMAT_BINARY 0x00000004
#define LINEADDRCAPFLAGS_FWDNUMRINGS 0x00000001
#define LINEADDRCAPFLAGS_PICKUPGROUPID 0x00000002
#define LINEADDRCAPFLAGS_SECURE 0x00000004
#define LINEADDRCAPFLAGS_BLOCKIDDEFAULT 0x00000008
#define LINEADDRCAPFLAGS_BLOCKIDOVERRIDE 0x00000010
#define LINEADDRCAPFLAGS_DIALED 0x00000020
#define LINEADDRCAPFLAGS_ORIGOFFHOOK 0x00000040
#define LINEADDRCAPFLAGS_DESTOFFHOOK 0x00000080
#define LINEADDRCAPFLAGS_FWDCONSULT 0x00000100
#define LINEADDRCAPFLAGS_SETUPCONFNULL 0x00000200
#define LINEADDRCAPFLAGS_AUTORECONNECT 0x00000400
#define LINEADDRCAPFLAGS_COMPLETIONID 0x00000800
#define LINEADDRCAPFLAGS_TRANSFERHELD 0x00001000
#define LINEADDRCAPFLAGS_TRANSFERMAKE 0x00002000
#define LINEADDRCAPFLAGS_CONFERENCEHELD 0x00004000
#define LINEADDRCAPFLAGS_CONFERENCEMAKE 0x00008000
#define LINEADDRCAPFLAGS_PARTIALDIAL 0x00010000
#define LINEADDRCAPFLAGS_FWDSTATUSVALID 0x00020000
#define LINEADDRCAPFLAGS_FWDINTEXTADDR 0x00040000
#define LINEADDRCAPFLAGS_FWDBUSYNAADDR 0x00080000
#define LINEADDRCAPFLAGS_ACCEPTTOALERT 0x00100000
#define LINEADDRCAPFLAGS_CONFDROP 0x00200000
#define LINEADDRCAPFLAGS_PICKUPCALLWAIT 0x00400000
#define LINEADDRESSMODE_ADDRESSID 0x00000001
#define LINEADDRESSMODE_DIALABLEADDR 0x00000002
#define LINEADDRESSSHARING_PRIVATE 0x00000001
#define LINEADDRESSSHARING_BRIDGEDEXCL 0x00000002
#define LINEADDRESSSHARING_BRIDGEDNEW 0x00000004
#define LINEADDRESSSHARING_BRIDGEDSHARED 0x00000008
#define LINEADDRESSSHARING_MONITORED 0x00000010
#define LINEADDRESSSTATE_OTHER 0x00000001
#define LINEADDRESSSTATE_DEVSPECIFIC 0x00000002
#define LINEADDRESSSTATE_INUSEZERO 0x00000004
#define LINEADDRESSSTATE_INUSEONE 0x00000008
#define LINEADDRESSSTATE_INUSEMANY 0x00000010
#define LINEADDRESSSTATE_NUMCALLS 0x00000020
#define LINEADDRESSSTATE_FORWARD 0x00000040
#define LINEADDRESSSTATE_TERMINALS 0x00000080
#define LINEADDRESSSTATE_CAPSCHANGE 0x00000100
#define LINEADDRFEATURE_FORWARD 0x00000001
#define LINEADDRFEATURE_MAKECALL 0x00000002
#define LINEADDRFEATURE_PICKUP 0x00000004
#define LINEADDRFEATURE_SETMEDIACONTROL 0x00000008
#define LINEADDRFEATURE_SETTERMINAL 0x00000010
#define LINEADDRFEATURE_SETUPCONF 0x00000020
#define LINEADDRFEATURE_UNCOMPLETECALL 0x00000040
#define LINEADDRFEATURE_UNPARK 0x00000080
#define LINEANSWERMODE_NONE 0x00000001
#define LINEANSWERMODE_DROP 0x00000002
#define LINEANSWERMODE_HOLD 0x00000004
#define LINEBEARERMODE_VOICE 0x00000001
#define LINEBEARERMODE_SPEECH 0x00000002
#define LINEBEARERMODE_MULTIUSE 0x00000004
#define LINEBEARERMODE_DATA 0x00000008
#define LINEBEARERMODE_ALTSPEECHDATA 0x00000010
#define LINEBEARERMODE_NONCALLSIGNALING 0x00000020
#define LINEBEARERMODE_PASSTHROUGH 0x00000040
#define LINEBUSYMODE_STATION 0x00000001
#define LINEBUSYMODE_TRUNK 0x00000002
#define LINEBUSYMODE_UNKNOWN 0x00000004
#define LINEBUSYMODE_UNAVAIL 0x00000008
#define LINECALLCOMPLCOND_BUSY 0x00000001
#define LINECALLCOMPLCOND_NOANSWER 0x00000002
#define LINECALLCOMPLMODE_CAMPON 0x00000001
#define LINECALLCOMPLMODE_CALLBACK 0x00000002
#define LINECALLCOMPLMODE_INTRUDE 0x00000004
#define LINECALLCOMPLMODE_MESSAGE 0x00000008
#define LINECALLFEATURE_ACCEPT 0x00000001
#define LINECALLFEATURE_ADDTOCONF 0x00000002
#define LINECALLFEATURE_ANSWER 0x00000004
#define LINECALLFEATURE_BLINDTRANSFER 0x00000008
#define LINECALLFEATURE_COMPLETECALL 0x00000010
#define LINECALLFEATURE_COMPLETETRANSF 0x00000020
#define LINECALLFEATURE_DIAL 0x00000040
#define LINECALLFEATURE_DROP 0x00000080
#define LINECALLFEATURE_GATHERDIGITS 0x00000100
#define LINECALLFEATURE_GENERATEDIGITS 0x00000200
#define LINECALLFEATURE_GENERATETONE 0x00000400
#define LINECALLFEATURE_HOLD 0x00000800
#define LINECALLFEATURE_MONITORDIGITS 0x00001000
#define LINECALLFEATURE_MONITORMEDIA 0x00002000
#define LINECALLFEATURE_MONITORTONES 0x00004000
#define LINECALLFEATURE_PARK 0x00008000
#define LINECALLFEATURE_PREPAREADDCONF 0x00010000
#define LINECALLFEATURE_REDIRECT 0x00020000
#define LINECALLFEATURE_REMOVEFROMCONF 0x00040000
#define LINECALLFEATURE_SECURECALL 0x00080000
#define LINECALLFEATURE_SENDUSERUSER 0x00100000
#define LINECALLFEATURE_SETCALLPARAMS 0x00200000
#define LINECALLFEATURE_SETMEDIACONTROL 0x00400000
#define LINECALLFEATURE_SETTERMINAL 0x00800000
#define LINECALLFEATURE_SETUPCONF 0x01000000
#define LINECALLFEATURE_SETUPTRANSFER 0x02000000
#define LINECALLFEATURE_SWAPHOLD 0x04000000
#define LINECALLFEATURE_UNHOLD 0x08000000
#define LINECALLFEATURE_RELEASEUSERUSERINFO 0x10000000
#define LINECALLINFOSTATE_OTHER 0x00000001
#define LINECALLINFOSTATE_DEVSPECIFIC 0x00000002
#define LINECALLINFOSTATE_BEARERMODE 0x00000004
#define LINECALLINFOSTATE_RATE 0x00000008
#define LINECALLINFOSTATE_MEDIAMODE 0x00000010
#define LINECALLINFOSTATE_APPSPECIFIC 0x00000020
#define LINECALLINFOSTATE_CALLID 0x00000040
#define LINECALLINFOSTATE_RELATEDCALLID 0x00000080
#define LINECALLINFOSTATE_ORIGIN 0x00000100
#define LINECALLINFOSTATE_REASON 0x00000200
#define LINECALLINFOSTATE_COMPLETIONID 0x00000400
#define LINECALLINFOSTATE_NUMOWNERINCR 0x00000800
#define LINECALLINFOSTATE_NUMOWNERDECR 0x00001000
#define LINECALLINFOSTATE_NUMMONITORS 0x00002000
#define LINECALLINFOSTATE_TRUNK 0x00004000
#define LINECALLINFOSTATE_CALLERID 0x00008000
#define LINECALLINFOSTATE_CALLEDID 0x00010000
#define LINECALLINFOSTATE_CONNECTEDID 0x00020000
#define LINECALLINFOSTATE_REDIRECTIONID 0x00040000
#define LINECALLINFOSTATE_REDIRECTINGID 0x00080000
#define LINECALLINFOSTATE_DISPLAY 0x00100000
#define LINECALLINFOSTATE_USERUSERINFO 0x00200000
#define LINECALLINFOSTATE_HIGHLEVELCOMP 0x00400000
#define LINECALLINFOSTATE_LOWLEVELCOMP 0x00800000
#define LINECALLINFOSTATE_CHARGINGINFO 0x01000000
#define LINECALLINFOSTATE_TERMINAL 0x02000000
#define LINECALLINFOSTATE_DIALPARAMS 0x04000000
#define LINECALLINFOSTATE_MONITORMODES 0x08000000
#define LINECALLORIGIN_OUTBOUND 0x00000001
#define LINECALLORIGIN_INTERNAL 0x00000002
#define LINECALLORIGIN_EXTERNAL 0x00000004
#define LINECALLORIGIN_UNKNOWN 0x00000010
#define LINECALLORIGIN_UNAVAIL 0x00000020
#define LINECALLORIGIN_CONFERENCE 0x00000040
#define LINECALLORIGIN_INBOUND 0x00000080
#define LINECALLPARAMFLAGS_SECURE 0x00000001
#define LINECALLPARAMFLAGS_IDLE 0x00000002
#define LINECALLPARAMFLAGS_BLOCKID 0x00000004
#define LINECALLPARAMFLAGS_ORIGOFFHOOK 0x00000008
#define LINECALLPARAMFLAGS_DESTOFFHOOK 0x00000010
#define LINECALLPARTYID_BLOCKED 0x00000001
#define LINECALLPARTYID_OUTOFAREA 0x00000002
#define LINECALLPARTYID_NAME 0x00000004
#define LINECALLPARTYID_ADDRESS 0x00000008
#define LINECALLPARTYID_PARTIAL 0x00000010
#define LINECALLPARTYID_UNKNOWN 0x00000020
#define LINECALLPARTYID_UNAVAIL 0x00000040
#define LINECALLPRIVILEGE_NONE 0x00000001
#define LINECALLPRIVILEGE_MONITOR 0x00000002
#define LINECALLPRIVILEGE_OWNER 0x00000004
#define LINECALLREASON_DIRECT 0x00000001
#define LINECALLREASON_FWDBUSY 0x00000002
#define LINECALLREASON_FWDNOANSWER 0x00000004
#define LINECALLREASON_FWDUNCOND 0x00000008
#define LINECALLREASON_PICKUP 0x00000010
#define LINECALLREASON_UNPARK 0x00000020
#define LINECALLREASON_REDIRECT 0x00000040
#define LINECALLREASON_CALLCOMPLETION 0x00000080
#define LINECALLREASON_TRANSFER 0x00000100
#define LINECALLREASON_REMINDER 0x00000200
#define LINECALLREASON_UNKNOWN 0x00000400
#define LINECALLREASON_UNAVAIL 0x00000800
#define LINECALLREASON_INTRUDE 0x00001000
#define LINECALLREASON_PARKED 0x00002000
#define LINECALLSELECT_LINE 0x00000001
#define LINECALLSELECT_ADDRESS 0x00000002
#define LINECALLSELECT_CALL 0x00000004
#define LINECALLSTATE_IDLE 0x00000001
#define LINECALLSTATE_OFFERING 0x00000002
#define LINECALLSTATE_ACCEPTED 0x00000004
#define LINECALLSTATE_DIALTONE 0x00000008
#define LINECALLSTATE_DIALING 0x00000010
#define LINECALLSTATE_RINGBACK 0x00000020
#define LINECALLSTATE_BUSY 0x00000040
#define LINECALLSTATE_SPECIALINFO 0x00000080
#define LINECALLSTATE_CONNECTED 0x00000100
#define LINECALLSTATE_PROCEEDING 0x00000200
#define LINECALLSTATE_ONHOLD 0x00000400
#define LINECALLSTATE_CONFERENCED 0x00000800
#define LINECALLSTATE_ONHOLDPENDCONF 0x00001000
#define LINECALLSTATE_ONHOLDPENDTRANSFER 0x00002000
#define LINECALLSTATE_DISCONNECTED 0x00004000
#define LINECALLSTATE_UNKNOWN 0x00008000
#define LINECONNECTEDMODE_ACTIVE 0x00000001
#define LINECONNECTEDMODE_INACTIVE 0x00000002
#define LINEOFFERINGMODE_ACTIVE 0x00000001
#define LINEOFFERINGMODE_INACTIVE 0x00000002
#define LINEDEVCAPFLAGS_CROSSADDRCONF 0x00000001
#define LINEDEVCAPFLAGS_HIGHLEVCOMP 0x00000002
#define LINEDEVCAPFLAGS_LOWLEVCOMP 0x00000004
#define LINEDEVCAPFLAGS_MEDIACONTROL 0x00000008
#define LINEDEVCAPFLAGS_MULTIPLEADDR 0x00000010
#define LINEDEVCAPFLAGS_CLOSEDROP 0x00000020
#define LINEDEVCAPFLAGS_DIALBILLING 0x00000040
#define LINEDEVCAPFLAGS_DIALQUIET 0x00000080
#define LINEDEVCAPFLAGS_DIALDIALTONE 0x00000100
#define LINEDEVSTATE_OTHER 0x00000001
#define LINEDEVSTATE_RINGING 0x00000002
#define LINEDEVSTATE_CONNECTED 0x00000004
#define LINEDEVSTATE_DISCONNECTED 0x00000008
#define LINEDEVSTATE_MSGWAITON 0x00000010
#define LINEDEVSTATE_MSGWAITOFF 0x00000020
#define LINEDEVSTATE_INSERVICE 0x00000040
#define LINEDEVSTATE_OUTOFSERVICE 0x00000080
#define LINEDEVSTATE_MAINTENANCE 0x00000100
#define LINEDEVSTATE_OPEN 0x00000200
#define LINEDEVSTATE_CLOSE 0x00000400
#define LINEDEVSTATE_NUMCALLS 0x00000800
#define LINEDEVSTATE_NUMCOMPLETIONS 0x00001000
#define LINEDEVSTATE_TERMINALS 0x00002000
#define LINEDEVSTATE_ROAMMODE 0x00004000
#define LINEDEVSTATE_BATTERY 0x00008000
#define LINEDEVSTATE_SIGNAL 0x00010000
#define LINEDEVSTATE_DEVSPECIFIC 0x00020000
#define LINEDEVSTATE_REINIT 0x00040000
#define LINEDEVSTATE_LOCK 0x00080000
#define LINEDEVSTATE_CAPSCHANGE 0x00100000
#define LINEDEVSTATE_CONFIGCHANGE 0x00200000
#define LINEDEVSTATE_TRANSLATECHANGE 0x00400000
#define LINEDEVSTATE_COMPLCANCEL 0x00800000
#define LINEDEVSTATE_REMOVED 0x01000000
#define LINEDEVSTATUSFLAGS_CONNECTED 0x00000001
#define LINEDEVSTATUSFLAGS_MSGWAIT 0x00000002
#define LINEDEVSTATUSFLAGS_INSERVICE 0x00000004
#define LINEDEVSTATUSFLAGS_LOCKED 0x00000008
#define LINEDIALTONEMODE_NORMAL 0x00000001
#define LINEDIALTONEMODE_SPECIAL 0x00000002
#define LINEDIALTONEMODE_INTERNAL 0x00000004
#define LINEDIALTONEMODE_EXTERNAL 0x00000008
#define LINEDIALTONEMODE_UNKNOWN 0x00000010
#define LINEDIALTONEMODE_UNAVAIL 0x00000020
#define LINEDIGITMODE_PULSE 0x00000001
#define LINEDIGITMODE_DTMF 0x00000002
#define LINEDIGITMODE_DTMFEND 0x00000004
#define LINEDISCONNECTMODE_NORMAL 0x00000001
#define LINEDISCONNECTMODE_UNKNOWN 0x00000002
#define LINEDISCONNECTMODE_REJECT 0x00000004
#define LINEDISCONNECTMODE_PICKUP 0x00000008
#define LINEDISCONNECTMODE_FORWARDED 0x00000010
#define LINEDISCONNECTMODE_BUSY 0x00000020
#define LINEDISCONNECTMODE_NOANSWER 0x00000040
#define LINEDISCONNECTMODE_BADADDRESS 0x00000080
#define LINEDISCONNECTMODE_UNREACHABLE 0x00000100
#define LINEDISCONNECTMODE_CONGESTION 0x00000200
#define LINEDISCONNECTMODE_INCOMPATIBLE 0x00000400
#define LINEDISCONNECTMODE_UNAVAIL 0x00000800
#define LINEDISCONNECTMODE_NODIALTONE 0x00001000
#define LINEERR_ALLOCATED 0x80000001
#define LINEERR_BADDEVICEID 0x80000002
#define LINEERR_BEARERMODEUNAVAIL 0x80000003
#define LINEERR_CALLUNAVAIL 0x80000005
#define LINEERR_COMPLETIONOVERRUN 0x80000006
#define LINEERR_CONFERENCEFULL 0x80000007
#define LINEERR_DIALBILLING 0x80000008
#define LINEERR_DIALDIALTONE 0x80000009
#define LINEERR_DIALPROMPT 0x8000000A
#define LINEERR_DIALQUIET 0x8000000B
#define LINEERR_INCOMPATIBLEAPIVERSION 0x8000000C
#define LINEERR_INCOMPATIBLEEXTVERSION 0x8000000D
#define LINEERR_INIFILECORRUPT 0x8000000E
#define LINEERR_INUSE 0x8000000F
#define LINEERR_INVALADDRESS 0x80000010
#define LINEERR_INVALADDRESSID 0x80000011
#define LINEERR_INVALADDRESSMODE 0x80000012
#define LINEERR_INVALADDRESSSTATE 0x80000013
#define LINEERR_INVALAPPHANDLE 0x80000014
#define LINEERR_INVALAPPNAME 0x80000015
#define LINEERR_INVALBEARERMODE 0x80000016
#define LINEERR_INVALCALLCOMPLMODE 0x80000017
#define LINEERR_INVALCALLHANDLE 0x80000018
#define LINEERR_INVALCALLPARAMS 0x80000019
#define LINEERR_INVALCALLPRIVILEGE 0x8000001A
#define LINEERR_INVALCALLSELECT 0x8000001B
#define LINEERR_INVALCALLSTATE 0x8000001C
#define LINEERR_INVALCALLSTATELIST 0x8000001D
#define LINEERR_INVALCARD 0x8000001E
#define LINEERR_INVALCOMPLETIONID 0x8000001F
#define LINEERR_INVALCONFCALLHANDLE 0x80000020
#define LINEERR_INVALCONSULTCALLHANDLE 0x80000021
#define LINEERR_INVALCOUNTRYCODE 0x80000022
#define LINEERR_INVALDEVICECLASS 0x80000023
#define LINEERR_INVALDEVICEHANDLE 0x80000024
#define LINEERR_INVALDIALPARAMS 0x80000025
#define LINEERR_INVALDIGITLIST 0x80000026
#define LINEERR_INVALDIGITMODE 0x80000027
#define LINEERR_INVALDIGITS 0x80000028
#define LINEERR_INVALEXTVERSION 0x80000029
#define LINEERR_INVALGROUPID 0x8000002A
#define LINEERR_INVALLINEHANDLE 0x8000002B
#define LINEERR_INVALLINESTATE 0x8000002C
#define LINEERR_INVALLOCATION 0x8000002D
#define LINEERR_INVALMEDIALIST 0x8000002E
#define LINEERR_INVALMEDIAMODE 0x8000002F
#define LINEERR_INVALMESSAGEID 0x80000030
#define LINEERR_INVALPARAM 0x80000032
#define LINEERR_INVALPARKID 0x80000033
#define LINEERR_INVALPARKMODE 0x80000034
#define LINEERR_INVALPOINTER 0x80000035
#define LINEERR_INVALPRIVSELECT 0x80000036
#define LINEERR_INVALRATE 0x80000037
#define LINEERR_INVALREQUESTMODE 0x80000038
#define LINEERR_INVALTERMINALID 0x80000039
#define LINEERR_INVALTERMINALMODE 0x8000003A
#define LINEERR_INVALTIMEOUT 0x8000003B
#define LINEERR_INVALTONE 0x8000003C
#define LINEERR_INVALTONELIST 0x8000003D
#define LINEERR_INVALTONEMODE 0x8000003E
#define LINEERR_INVALTRANSFERMODE 0x8000003F
#define LINEERR_LINEMAPPERFAILED 0x80000040
#define LINEERR_NOCONFERENCE 0x80000041
#define LINEERR_NODEVICE 0x80000042
#define LINEERR_NODRIVER 0x80000043
#define LINEERR_NOMEM 0x80000044
#define LINEERR_NOREQUEST 0x80000045
#define LINEERR_NOTOWNER 0x80000046
#define LINEERR_NOTREGISTERED 0x80000047
#define LINEERR_OPERATIONFAILED 0x80000048
#define LINEERR_OPERATIONUNAVAIL 0x80000049
#define LINEERR_RATEUNAVAIL 0x8000004A
#define LINEERR_RESOURCEUNAVAIL 0x8000004B
#define LINEERR_REQUESTOVERRUN 0x8000004C
#define LINEERR_STRUCTURETOOSMALL 0x8000004D
#define LINEERR_TARGETNOTFOUND 0x8000004E
#define LINEERR_TARGETSELF 0x8000004F
#define LINEERR_UNINITIALIZED 0x80000050
#define LINEERR_USERUSERINFOTOOBIG 0x80000051
#define LINEERR_REINIT 0x80000052
#define LINEERR_ADDRESSBLOCKED 0x80000053
#define LINEERR_BILLINGREJECTED 0x80000054
#define LINEERR_INVALFEATURE 0x80000055
#define LINEERR_NOMULTIPLEINSTANCE 0x80000056
#define LINEFEATURE_DEVSPECIFIC 0x00000001
#define LINEFEATURE_DEVSPECIFICFEAT 0x00000002
#define LINEFEATURE_FORWARD 0x00000004
#define LINEFEATURE_MAKECALL 0x00000008
#define LINEFEATURE_SETMEDIACONTROL 0x00000010
#define LINEFEATURE_SETTERMINAL 0x00000020
#define LINEFORWARDMODE_UNCOND 0x00000001
#define LINEFORWARDMODE_UNCONDINTERNAL 0x00000002
#define LINEFORWARDMODE_UNCONDEXTERNAL 0x00000004
#define LINEFORWARDMODE_UNCONDSPECIFIC 0x00000008
#define LINEFORWARDMODE_BUSY 0x00000010
#define LINEFORWARDMODE_BUSYINTERNAL 0x00000020
#define LINEFORWARDMODE_BUSYEXTERNAL 0x00000040
#define LINEFORWARDMODE_BUSYSPECIFIC 0x00000080
#define LINEFORWARDMODE_NOANSW 0x00000100
#define LINEFORWARDMODE_NOANSWINTERNAL 0x00000200
#define LINEFORWARDMODE_NOANSWEXTERNAL 0x00000400
#define LINEFORWARDMODE_NOANSWSPECIFIC 0x00000800
#define LINEFORWARDMODE_BUSYNA 0x00001000
#define LINEFORWARDMODE_BUSYNAINTERNAL 0x00002000
#define LINEFORWARDMODE_BUSYNAEXTERNAL 0x00004000
#define LINEFORWARDMODE_BUSYNASPECIFIC 0x00008000
#define LINEFORWARDMODE_UNKNOWN 0x00010000
#define LINEFORWARDMODE_UNAVAIL 0x00020000
#define LINEGATHERTERM_BUFFERFULL 0x00000001
#define LINEGATHERTERM_TERMDIGIT 0x00000002
#define LINEGATHERTERM_FIRSTTIMEOUT 0x00000004
#define LINEGATHERTERM_INTERTIMEOUT 0x00000008
#define LINEGATHERTERM_CANCEL 0x00000010
#define LINEGENERATETERM_DONE 0x00000001
#define LINEGENERATETERM_CANCEL 0x00000002
#define LINEMEDIACONTROL_NONE 0x00000001
#define LINEMEDIACONTROL_START 0x00000002
#define LINEMEDIACONTROL_RESET 0x00000004
#define LINEMEDIACONTROL_PAUSE 0x00000008
#define LINEMEDIACONTROL_RESUME 0x00000010
#define LINEMEDIACONTROL_RATEUP 0x00000020
#define LINEMEDIACONTROL_RATEDOWN 0x00000040
#define LINEMEDIACONTROL_RATENORMAL 0x00000080
#define LINEMEDIACONTROL_VOLUMEUP 0x00000100
#define LINEMEDIACONTROL_VOLUMEDOWN 0x00000200
#define LINEMEDIACONTROL_VOLUMENORMAL 0x00000400
#define LINEMEDIAMODE_UNKNOWN 0x00000002
#define LINEMEDIAMODE_INTERACTIVEVOICE 0x00000004
#define LINEMEDIAMODE_AUTOMATEDVOICE 0x00000008
#define LINEMEDIAMODE_DATAMODEM 0x00000010
#define LINEMEDIAMODE_G3FAX 0x00000020
#define LINEMEDIAMODE_TDD 0x00000040
#define LINEMEDIAMODE_G4FAX 0x00000080
#define LINEMEDIAMODE_DIGITALDATA 0x00000100
#define LINEMEDIAMODE_TELETEX 0x00000200
#define LINEMEDIAMODE_VIDEOTEX 0x00000400
#define LINEMEDIAMODE_TELEX 0x00000800
#define LINEMEDIAMODE_MIXED 0x00001000
#define LINEMEDIAMODE_ADSI 0x00002000
#define LINEMEDIAMODE_VOICEVIEW 0x00004000
#define LAST_LINEMEDIAMODE 0x00004000
#define LINEPARKMODE_DIRECTED 0x00000001
#define LINEPARKMODE_NONDIRECTED 0x00000002
#define LINEREMOVEFROMCONF_NONE 0x00000001
#define LINEREMOVEFROMCONF_LAST 0x00000002
#define LINEREMOVEFROMCONF_ANY 0x00000003
#define LINEREQUESTMODE_MAKECALL 0x00000001
#define LINEREQUESTMODE_MEDIACALL 0x00000002
#define LINEREQUESTMODE_DROP 0x00000004
#define LAST_LINEREQUESTMODE LINEREQUESTMODE_MEDIACALL
#define LINEROAMMODE_UNKNOWN 0x00000001
#define LINEROAMMODE_UNAVAIL 0x00000002
#define LINEROAMMODE_HOME 0x00000004
#define LINEROAMMODE_ROAMA 0x00000008
#define LINEROAMMODE_ROAMB 0x00000010
#define LINESPECIALINFO_NOCIRCUIT 0x00000001
#define LINESPECIALINFO_CUSTIRREG 0x00000002
#define LINESPECIALINFO_REORDER 0x00000004
#define LINESPECIALINFO_UNKNOWN 0x00000008
#define LINESPECIALINFO_UNAVAIL 0x00000010
#define LINETERMDEV_PHONE 0x00000001
#define LINETERMDEV_HEADSET 0x00000002
#define LINETERMDEV_SPEAKER 0x00000004
#define LINETERMMODE_BUTTONS 0x00000001
#define LINETERMMODE_LAMPS 0x00000002
#define LINETERMMODE_DISPLAY 0x00000004
#define LINETERMMODE_RINGER 0x00000008
#define LINETERMMODE_HOOKSWITCH 0x00000010
#define LINETERMMODE_MEDIATOLINE 0x00000020
#define LINETERMMODE_MEDIAFROMLINE 0x00000040
#define LINETERMMODE_MEDIABIDIRECT 0x00000080
#define LINETERMSHARING_PRIVATE 0x00000001
#define LINETERMSHARING_SHAREDEXCL 0x00000002
#define LINETERMSHARING_SHAREDCONF 0x00000004
#define LINETONEMODE_CUSTOM 0x00000001
#define LINETONEMODE_RINGBACK 0x00000002
#define LINETONEMODE_BUSY 0x00000004
#define LINETONEMODE_BEEP 0x00000008
#define LINETONEMODE_BILLING 0x00000010
#define LINETRANSFERMODE_TRANSFER 0x00000001
#define LINETRANSFERMODE_CONFERENCE 0x00000002
#define LINETOLLLISTOPTION_ADD 0x00000001
#define LINETOLLLISTOPTION_REMOVE 0x00000002
#define LINETRANSLATEOPTION_CARDOVERRIDE 0x00000001
#define LINETRANSLATEOPTION_CANCELCALLWAITING 0x00000002
#define LINETRANSLATEOPTION_FORCELOCAL 0x00000004
#define LINETRANSLATEOPTION_FORCELD 0x00000008
#define LINETRANSLATERESULT_CANONICAL 0x00000001
#define LINETRANSLATERESULT_INTERNATIONAL 0x00000002
#define LINETRANSLATERESULT_LONGDISTANCE 0x00000004
#define LINETRANSLATERESULT_LOCAL 0x00000008
#define LINETRANSLATERESULT_INTOLLLIST 0x00000010
#define LINETRANSLATERESULT_NOTINTOLLLIST 0x00000020
#define LINETRANSLATERESULT_DIALBILLING 0x00000040
#define LINETRANSLATERESULT_DIALQUIET 0x00000080
#define LINETRANSLATERESULT_DIALDIALTONE 0x00000100
#define LINETRANSLATERESULT_DIALPROMPT 0x00000200
#define LINELOCATIONOPTION_PULSEDIAL 0x00000001
#define LINECARDOPTION_PREDEFINED 0x00000001
#define LINECARDOPTION_HIDDEN 0x00000002
#define INVALID_HANDLE_VALUE PTR (_CAST, 0xFFFFFFFF)
#define INVALID_FILE_SIZE DWORD (_CAST, 0xFFFFFFFF)
#define FILE_BEGIN 0
#define FILE_CURRENT 1
#define FILE_END 2
#define TIME_ZONE_ID_INVALID DWORD (_CAST, 0xFFFFFFFF)
#define WAIT_FAILED DWORD (_CAST, 0xFFFFFFFF)
#define STATUS_WAIT_0 0x00000000L
#define WAIT_OBJECT_0 STATUS_WAIT_0 + 0
#define STATUS_ABANDONED_WAIT_0 0x00000080L
#define WAIT_ABANDONED (STATUS_ABANDONED_WAIT_0 + 0 )
#define WAIT_ABANDONED_0 (STATUS_ABANDONED_WAIT_0 + 0 )
#define STATUS_TIMEOUT DWORD (_CAST, 0x00000102L)
#define WAIT_TIMEOUT STATUS_TIMEOUT
#define STATUS_USER_APC DWORD (_CAST, 0x000000C0)
#define WAIT_IO_COMPLETION STATUS_USER_APC
#define STATUS_PENDING DWORD (_CAST, 0x00000103L)
#define STILL_ACTIVE STATUS_PENDING
#define STATUS_ACCESS_VIOLATION DWORD (_CAST, 0xC0000005L)
#define EXCEPTION_ACCESS_VIOLATION STATUS_ACCESS_VIOLATION
#define STATUS_DATATYPE_MISALIGNMENT DWORD (_CAST, 0x80000002L)
#define EXCEPTION_DATATYPE_MISALIGNMENT STATUS_DATATYPE_MISALIGNMENT
#define STATUS_BREAKPOINT DWORD (_CAST, 0x80000003L)
#define EXCEPTION_BREAKPOINT STATUS_BREAKPOINT
#define STATUS_SINGLE_STEP DWORD (_CAST, 0x80000004L)
#define EXCEPTION_SINGLE_STEP STATUS_SINGLE_STEP
#define STATUS_ARRAY_BOUNDS_EXCEEDED DWORD (_CAST, 0xC000008CL)
#define EXCEPTION_ARRAY_BOUNDS_EXCEEDED STATUS_ARRAY_BOUNDS_EXCEEDED
#define STATUS_FLOAT_DENORMAL_OPERAND DWORD (_CAST, 0xC000008DL)
#define EXCEPTION_FLT_DENORMAL_OPERAND STATUS_FLOAT_DENORMAL_OPERAND
#define STATUS_FLOAT_DIVIDE_BY_ZERO DWORD (_CAST, 0xC000008EL)
#define EXCEPTION_FLT_DIVIDE_BY_ZERO STATUS_FLOAT_DIVIDE_BY_ZERO
#define STATUS_FLOAT_INEXACT_RESULT DWORD (_CAST, 0xC000008FL)
#define EXCEPTION_FLT_INEXACT_RESULT STATUS_FLOAT_INEXACT_RESULT
#define STATUS_FLOAT_INVALID_OPERATION DWORD (_CAST, 0xC0000090L)
#define EXCEPTION_FLT_INVALID_OPERATION STATUS_FLOAT_INVALID_OPERATION
#define STATUS_FLOAT_OVERFLOW DWORD (_CAST, 0xC0000091L)
#define EXCEPTION_FLT_OVERFLOW STATUS_FLOAT_OVERFLOW
#define STATUS_FLOAT_STACK_CHECK DWORD (_CAST, 0xC0000092L)
#define EXCEPTION_FLT_STACK_CHECK STATUS_FLOAT_STACK_CHECK
#define STATUS_FLOAT_UNDERFLOW DWORD (_CAST, 0xC0000093L)
#define EXCEPTION_FLT_UNDERFLOW STATUS_FLOAT_UNDERFLOW
#define STATUS_INTEGER_DIVIDE_BY_ZERO DWORD (_CAST, 0xC0000094L)
#define EXCEPTION_INT_DIVIDE_BY_ZERO STATUS_INTEGER_DIVIDE_BY_ZERO
#define STATUS_INTEGER_OVERFLOW DWORD (_CAST, 0xC0000095L)
#define EXCEPTION_INT_OVERFLOW STATUS_INTEGER_OVERFLOW
#define STATUS_PRIVILEGED_INSTRUCTION DWORD (_CAST, 0xC0000096L)
#define EXCEPTION_PRIV_INSTRUCTION STATUS_PRIVILEGED_INSTRUCTION
#define STATUS_IN_PAGE_ERROR DWORD (_CAST, 0xC0000006L)
#define EXCEPTION_IN_PAGE_ERROR STATUS_IN_PAGE_ERROR
#define STATUS_ILLEGAL_INSTRUCTION DWORD (_CAST, 0xC000001DL)
#define EXCEPTION_ILLEGAL_INSTRUCTION STATUS_ILLEGAL_INSTRUCTION
#define STATUS_NONCONTINUABLE_EXCEPTION DWORD (_CAST, 0xC0000025L)
#define EXCEPTION_NONCONTINUABLE_EXCEPTION STATUS_NONCONTINUABLE_EXCEPTION
#define STATUS_STACK_OVERFLOW DWORD (_CAST, 0xC00000FDL)
#define EXCEPTION_STACK_OVERFLOW STATUS_STACK_OVERFLOW
#define STATUS_INVALID_DISPOSITION DWORD (_CAST, 0xC0000026L)
#define EXCEPTION_INVALID_DISPOSITION STATUS_INVALID_DISPOSITION
#define STATUS_GUARD_PAGE_VIOLATION DWORD (_CAST, 0x80000001L)
#define EXCEPTION_GUARD_PAGE STATUS_GUARD_PAGE_VIOLATION
#define STATUS_CONTROL_C_EXIT DWORD (_CAST, 0xC000013AL)
#define CONTROL_C_EXIT STATUS_CONTROL_C_EXIT
#define FILE_FLAG_WRITE_THROUGH 0x80000000
#define FILE_FLAG_OVERLAPPED 0x40000000
#define FILE_FLAG_NO_BUFFERING 0x20000000
#define FILE_FLAG_RANDOM_ACCESS 0x10000000
#define FILE_FLAG_SEQUENTIAL_SCAN 0x08000000
#define FILE_FLAG_DELETE_ON_CLOSE 0x04000000
#define FILE_FLAG_BACKUP_SEMANTICS 0x02000000
#define FILE_FLAG_POSIX_SEMANTICS 0x01000000
#define CREATE_NEW 1
#define CREATE_ALWAYS 2
#define OPEN_EXISTING 3
#define OPEN_ALWAYS 4
#define TRUNCATE_EXISTING 5
#define PIPE_ACCESS_INBOUND 0x00000001
#define PIPE_ACCESS_OUTBOUND 0x00000002
#define PIPE_ACCESS_DUPLEX 0x00000003
#define PIPE_CLIENT_END 0x00000000
#define PIPE_SERVER_END 0x00000001
#define PIPE_WAIT 0x00000000
#define PIPE_NOWAIT 0x00000001
#define PIPE_READMODE_BYTE 0x00000000
#define PIPE_READMODE_MESSAGE 0x00000002
#define PIPE_TYPE_MESSAGE 0x00000004
#define PIPE_UNLIMITED_INSTANCES 255
#define SECURITY_SQOS_PRESENT 0x00100000
#define SECURITY_VALID_SQOS_FLAGS 0x001F0000
#define MUTANT_QUERY_STATE 0x0001
#define MUTEX_MODIFY_STATE MUTANT_QUERY_STATE
#define MUTANT_ALL_ACCESS 0x001F0001
#define MUTEX_ALL_ACCESS MUTANT_ALL_ACCESS
#define COMMPROP_INITIALIZED DWORD(_CAST, 0xE73CF52E)
#define DTR_CONTROL_DISABLE 0x00
#define DTR_CONTROL_ENABLE 0x01
#define DTR_CONTROL_HANDSHAKE 0x02
#define RTS_CONTROL_DISABLE 0x00
#define RTS_CONTROL_ENABLE 0x01
#define RTS_CONTROL_HANDSHAKE 0x02
#define RTS_CONTROL_TOGGLE 0x03
#define GMEM_FIXED 0x0000
#define GMEM_MOVEABLE 0x0002
#define GMEM_NOCOMPACT 0x0010
#define GMEM_NODISCARD 0x0020
#define GMEM_ZEROINIT 0x0040
#define GMEM_MODIFY 0x0080
#define GMEM_DISCARDABLE 0x0100
#define GMEM_NOT_BANKED 0x1000
#define GMEM_SHARE 0x2000
#define GMEM_DDESHARE 0x2000
#define GMEM_NOTIFY 0x4000
#define GMEM_LOWER GMEM_NOT_BANKED
#define GMEM_VALID_FLAGS 0x7F72
#define GMEM_INVALID_HANDLE 0x8000
#define GHND 0x0042
#define GPTR 0x0040
#define GMEM_DISCARDED 0x4000
#define GMEM_LOCKCOUNT 0x00FF
#define LMEM_FIXED 0x0000
#define LMEM_MOVEABLE 0x0002
#define LMEM_NOCOMPACT 0x0010
#define LMEM_NODISCARD 0x0020
#define LMEM_ZEROINIT 0x0040
#define LMEM_MODIFY 0x0080
#define LMEM_DISCARDABLE 0x0F00
#define LMEM_VALID_FLAGS 0x0F72
#define LMEM_INVALID_HANDLE 0x8000
#define LHND 0x0042
#define LPTR 0x0040
#define NONZEROLHND (LMEM_MOVEABLE)
#define NONZEROLPTR (LMEM_FIXED)
#define LMEM_DISCARDED 0x4000
#define LMEM_LOCKCOUNT 0x00FF
#define DEBUG_PROCESS 0x00000001
#define DEBUG_ONLY_THIS_PROCESS 0x00000002
#define CREATE_SUSPENDED 0x00000004
#define DETACHED_PROCESS 0x00000008
#define CREATE_NEW_CONSOLE 0x00000010
#define NORMAL_PRIORITY_CLASS 0x00000020
#define IDLE_PRIORITY_CLASS 0x00000040
#define HIGH_PRIORITY_CLASS 0x00000080
#define REALTIME_PRIORITY_CLASS 0x00000100
#define CREATE_NEW_PROCESS_GROUP 0x00000200
#define CREATE_UNICODE_ENVIRONMENT 0x00000400
#define CREATE_SEPARATE_WOW_VDM 0x00000800
#define CREATE_SHARED_WOW_VDM 0x00001000
#define CREATE_DEFAULT_ERROR_MODE 0x04000000
#define CREATE_NO_WINDOW 0x08000000
#define PROFILE_USER 0x10000000
#define PROFILE_KERNEL 0x20000000
#define PROFILE_SERVER 0x40000000
#define THREAD_BASE_PRIORITY_MIN -2
#define THREAD_PRIORITY_LOWEST THREAD_BASE_PRIORITY_MIN
#define THREAD_PRIORITY_BELOW_NORMAL (THREAD_PRIORITY_LOWEST+1)
#define THREAD_PRIORITY_NORMAL 0
#define THREAD_BASE_PRIORITY_MAX 2
#define THREAD_PRIORITY_HIGHEST THREAD_BASE_PRIORITY_MAX
#define THREAD_PRIORITY_ABOVE_NORMAL (THREAD_PRIORITY_HIGHEST-1)
#define MAXLONG 0x7fffffff
#define THREAD_PRIORITY_ERROR_RETURN (MAXLONG)
#define THREAD_BASE_PRIORITY_LOWRT 15
#define THREAD_PRIORITY_TIME_CRITICAL THREAD_BASE_PRIORITY_LOWRT
#define THREAD_BASE_PRIORITY_IDLE -15
#define THREAD_PRIORITY_IDLE THREAD_BASE_PRIORITY_IDLE
#define EXCEPTION_DEBUG_EVENT 1
#define CREATE_THREAD_DEBUG_EVENT 2
#define CREATE_PROCESS_DEBUG_EVENT 3
#define EXIT_THREAD_DEBUG_EVENT 4
#define EXIT_PROCESS_DEBUG_EVENT 5
#define LOAD_DLL_DEBUG_EVENT 6
#define UNLOAD_DLL_DEBUG_EVENT 7
#define OUTPUT_DEBUG_STRING_EVENT 8
#define RIP_EVENT 9
#define DRIVE_UNKNOWN 0
#define DRIVE_NO_ROOT_DIR 1
#define DRIVE_REMOVABLE 2
#define DRIVE_FIXED 3
#define DRIVE_REMOTE 4
#define DRIVE_CDROM 5
#define DRIVE_RAMDISK 6
#define FILE_TYPE_UNKNOWN 0x0000
#define FILE_TYPE_DISK 0x0001
#define FILE_TYPE_CHAR 0x0002
#define FILE_TYPE_PIPE 0x0003
#define FILE_TYPE_REMOTE 0x8000
#define STD_INPUT_HANDLE 0xFFFFFFF6
#define STD_OUTPUT_HANDLE 0xFFFFFFF5
#define STD_ERROR_HANDLE 0xFFFFFFF4
#define NOPARITY 0
#define ODDPARITY 1
#define EVENPARITY 2
#define MARKPARITY 3
#define SPACEPARITY 4
#define ONESTOPBIT 0
#define ONE5STOPBITS 1
#define TWOSTOPBITS 2
#define IGNORE 0
#define INFINITE DWORD(_CAST, 0xFFFFFFFF )
#define CBR_110 110
#define CBR_300 300
#define CBR_600 600
#define CBR_1200 1200
#define CBR_2400 2400
#define CBR_4800 4800
#define CBR_9600 9600
#define CBR_14400 14400
#define CBR_19200 19200
#define CBR_38400 38400
#define CBR_56000 56000
#define CBR_57600 57600
#define CBR_115200 115200
#define CBR_128000 128000
#define CBR_256000 256000
#define CBR_28800 28800
#define CE_RXOVER 0x0001
#define CE_OVERRUN 0x0002
#define CE_RXPARITY 0x0004
#define CE_FRAME 0x0008
#define CE_BREAK 0x0010
#define CE_TXFULL 0x0100
#define CE_PTO 0x0200
#define CE_IOE 0x0400
#define CE_DNS 0x0800
#define CE_OOP 0x1000
#define CE_MODE 0x8000
#define IE_BADID (-1)
#define IE_OPEN (-2)
#define IE_NOPEN (-3)
#define IE_MEMORY (-4)
#define IE_DEFAULT (-5)
#define IE_HARDWARE (-10)
#define IE_BYTESIZE (-11)
#define IE_BAUDRATE (-12)
#define EV_RXCHAR 0x0001
#define EV_RXFLAG 0x0002
#define EV_TXEMPTY 0x0004
#define EV_CTS 0x0008
#define EV_DSR 0x0010
#define EV_RLSD 0x0020
#define EV_BREAK 0x0040
#define EV_ERR 0x0080
#define EV_RING 0x0100
#define EV_PERR 0x0200
#define EV_RX80FULL 0x0400
#define EV_EVENT1 0x0800
#define EV_EVENT2 0x1000
#define SETXOFF 1
#define SETXON 2
#define SETRTS 3
#define CLRRTS 4
#define SETDTR 5
#define CLRDTR 6
#define RESETDEV 7
#define SETBREAK 8
#define CLRBREAK 9
#define PURGE_TXABORT 0x0001
#define PURGE_RXABORT 0x0002
#define PURGE_TXCLEAR 0x0004
#define PURGE_RXCLEAR 0x0008
#define LPTx 0x80
#define MS_CTS_ON DWORD (_CAST, 0x0010)
#define MS_DSR_ON DWORD (_CAST, 0x0020)
#define MS_RING_ON DWORD (_CAST, 0x0040)
#define MS_RLSD_ON DWORD (_CAST, 0x0080)
#define S_QUEUEEMPTY 0
#define S_THRESHOLD 1
#define S_ALLTHRESHOLD 2
#define S_NORMAL 0
#define S_LEGATO 1
#define S_STACCATO 2
#define S_PERIOD512 0
#define S_PERIOD1024 1
#define S_PERIOD2048 2
#define S_PERIODVOICE 3
#define S_WHITE512 4
#define S_WHITE1024 5
#define S_WHITE2048 6
#define S_WHITEVOICE 7
#define S_SERDVNA (-1)
#define S_SEROFM (-2)
#define S_SERMACT (-3)
#define S_SERQFUL (-4)
#define S_SERBDNT (-5)
#define S_SERDLN (-6)
#define S_SERDCC (-7)
#define S_SERDTP (-8)
#define S_SERDVL (-9)
#define S_SERDMD (-10)
#define S_SERDSH (-11)
#define S_SERDPT (-12)
#define S_SERDFQ (-13)
#define S_SERDDR (-14)
#define S_SERDSR (-15)
#define S_SERDST (-16)
#define NMPWAIT_WAIT_FOREVER 0xffffffff
#define NMPWAIT_NOWAIT 0x00000001
#define NMPWAIT_USE_DEFAULT_WAIT 0x00000000
#define FILE_CASE_PRESERVED_NAMES 0x00000002
#define FS_CASE_IS_PRESERVED FILE_CASE_PRESERVED_NAMES
#define FILE_CASE_SENSITIVE_SEARCH 0x00000001
#define FS_CASE_SENSITIVE FILE_CASE_SENSITIVE_SEARCH
#define FILE_UNICODE_ON_DISK 0x00000004
#define FS_UNICODE_STORED_ON_DISK FILE_UNICODE_ON_DISK
#define FILE_PERSISTENT_ACLS 0x00000008
#define FS_PERSISTENT_ACLS FILE_PERSISTENT_ACLS
#define FILE_VOLUME_IS_COMPRESSED 0x00008000
#define FS_VOL_IS_COMPRESSED FILE_VOLUME_IS_COMPRESSED
#define FILE_FILE_COMPRESSION 0x00000010
#define FS_FILE_COMPRESSION FILE_FILE_COMPRESSION
#define SECTION_QUERY 0x0001
#define FILE_MAP_COPY SECTION_QUERY
#define SECTION_MAP_WRITE 0x0002
#define FILE_MAP_WRITE SECTION_MAP_WRITE
#define SECTION_MAP_READ 0x0004
#define FILE_MAP_READ SECTION_MAP_READ
#define SECTION_ALL_ACCESS 0x000F001Fl
#define FILE_MAP_ALL_ACCESS SECTION_ALL_ACCESS
#define OF_READ 0x00000000
#define OF_WRITE 0x00000001
#define OF_READWRITE 0x00000002
#define OF_SHARE_COMPAT 0x00000000
#define OF_SHARE_EXCLUSIVE 0x00000010
#define OF_SHARE_DENY_WRITE 0x00000020
#define OF_SHARE_DENY_READ 0x00000030
#define OF_SHARE_DENY_NONE 0x00000040
#define OF_PARSE 0x00000100
#define OF_DELETE 0x00000200
#define OF_VERIFY 0x00000400
#define OF_CANCEL 0x00000800
#define OF_CREATE 0x00001000
#define OF_PROMPT 0x00002000
#define OF_EXIST 0x00004000
#define OF_REOPEN 0x00008000
#define OFS_MAXPATHNAME 128
#define MAXINTATOM 0xC000
#define PROCESS_HEAP_REGION 0x0001
#define PROCESS_HEAP_UNCOMMITTED_RANGE 0x0002
#define PROCESS_HEAP_ENTRY_BUSY 0x0004
#define PROCESS_HEAP_ENTRY_MOVEABLE 0x0010
#define PROCESS_HEAP_ENTRY_DDESHARE 0x0020
#define SCS_32BIT_BINARY 0
#define SCS_DOS_BINARY 1
#define SCS_WOW_BINARY 2
#define SCS_PIF_BINARY 3
#define SCS_POSIX_BINARY 4
#define SCS_OS216_BINARY 5
#define SEM_FAILCRITICALERRORS 0x0001
#define SEM_NOGPFAULTERRORBOX 0x0002
#define SEM_NOALIGNMENTFAULTEXCEPT 0x0004
#define SEM_NOOPENFILEERRORBOX 0x8000
#define LOCKFILE_FAIL_IMMEDIATELY 0x00000001
#define LOCKFILE_EXCLUSIVE_LOCK 0x00000002
#define HANDLE_FLAG_INHERIT 0x00000001
#define HANDLE_FLAG_PROTECT_FROM_CLOSE 0x00000002
#define HINSTANCE_ERROR 32
#define GET_TAPE_MEDIA_INFORMATION 0
#define GET_TAPE_DRIVE_INFORMATION 1
#define SET_TAPE_MEDIA_INFORMATION 0
#define SET_TAPE_DRIVE_INFORMATION 1
#define FORMAT_MESSAGE_ALLOCATE_BUFFER 0x00000100
#define FORMAT_MESSAGE_IGNORE_INSERTS 0x00000200
#define FORMAT_MESSAGE_FROM_STRING 0x00000400
#define FORMAT_MESSAGE_FROM_HMODULE 0x00000800
#define FORMAT_MESSAGE_FROM_SYSTEM 0x00001000
#define FORMAT_MESSAGE_ARGUMENT_ARRAY 0x00002000
#define FORMAT_MESSAGE_MAX_WIDTH_MASK 0x000000FF
#define TLS_OUT_OF_INDEXES DWORD(_CAST,0xFFFFFFFF)
#define BACKUP_INVALID 0x00000000
#define BACKUP_DATA 0x00000001
#define BACKUP_EA_DATA 0x00000002
#define BACKUP_SECURITY_DATA 0x00000003
#define BACKUP_ALTERNATE_DATA 0x00000004
#define BACKUP_LINK 0x00000005
#define BACKUP_PROPERTY_DATA 0x00000006
#define STREAM_NORMAL_ATTRIBUTE 0x00000000
#define STREAM_MODIFIED_WHEN_READ 0x00000001
#define STREAM_CONTAINS_SECURITY 0x00000002
#define STREAM_CONTAINS_PROPERTIES 0x00000004
#define STARTF_USESHOWWINDOW 0x00000001
#define STARTF_USESIZE 0x00000002
#define STARTF_USEPOSITION 0x00000004
#define STARTF_USECOUNTCHARS 0x00000008
#define STARTF_USEFILLATTRIBUTE 0x00000010
#define STARTF_RUNFULLSCREEN 0x00000020
#define STARTF_FORCEONFEEDBACK 0x00000040
#define STARTF_FORCEOFFFEEDBACK 0x00000080
#define STARTF_USESTDHANDLES 0x00000100
#define STARTF_USEHOTKEY 0x00000200
#define SHUTDOWN_NORETRY 0x00000001
#define DONT_RESOLVE_DLL_REFERENCES 0x00000001
#define LOAD_LIBRARY_AS_DATAFILE 0x00000002
#define LOAD_WITH_ALTERED_SEARCH_PATH 0x00000008
#define DDD_RAW_TARGET_PATH 0x00000001
#define DDD_REMOVE_DEFINITION 0x00000002
#define DDD_EXACT_MATCH_ON_REMOVE 0x00000004
#define MOVEFILE_REPLACE_EXISTING 0x00000001
#define MOVEFILE_COPY_ALLOWED 0x00000002
#define MOVEFILE_DELAY_UNTIL_REBOOT 0x00000004
#define MAX_COMPUTERNAME_LENGTH 15
#define LOGON32_LOGON_INTERACTIVE 2
#define LOGON32_LOGON_BATCH 4
#define LOGON32_LOGON_SERVICE 5
#define LOGON32_PROVIDER_DEFAULT 0
#define LOGON32_PROVIDER_WINNT35 1
#define VER_PLATFORM_WIN32s 0
#define VER_PLATFORM_WIN32_WINDOWS 1
#define VER_PLATFORM_WIN32_NT 2
#define TC_NORMAL 0
#define TC_HARDERR 1
#define TC_GP_TRAP 2
#define TC_SIGNAL 3
#define AC_LINE_OFFLINE 0x00
#define AC_LINE_ONLINE 0x01
#define AC_LINE_BACKUP_POWER 0x02
#define AC_LINE_UNKNOWN 0xFF
#define BATTERY_FLAG_HIGH 0x01
#define BATTERY_FLAG_LOW 0x02
#define BATTERY_FLAG_CRITICAL 0x04
#define BATTERY_FLAG_CHARGING 0x08
#define BATTERY_FLAG_NO_BATTERY 0x80
#define BATTERY_FLAG_UNKNOWN 0xFF
#define BATTERY_PERCENTAGE_UNKNOWN 0xFF
#define BATTERY_LIFE_UNKNOWN 0xFFFFFFFF
#define VER_NT_WORKSTATION 0x0000001
#define VER_NT_DOMAIN_CONTROLLER 0x0000002
#define VER_NT_SERVER 0x0000003
#define VER_SERVER_NT 0x80000000
#define VER_WORKSTATION_NT 0x40000000
#define VER_SUITE_SMALLBUSINESS 0x00000001
#define VER_SUITE_ENTERPRISE 0x00000002
#define VER_SUITE_BACKOFFICE 0x00000004
#define VER_SUITE_COMMUNICATIONS 0x00000008
#define VER_SUITE_TERMINAL 0x00000010
#define VER_SUITE_SMALLBUSINESS_RESTRICTED 0x00000020
#define VER_SUITE_EMBEDDEDNT 0x00000040
#define VER_SUITE_DATACENTER 0x00000080
#define VER_SUITE_SINGLEUSERTS 0x00000100
#define VER_SUITE_PERSONAL 0x00000200
#define VER_SUITE_BLADE 0x00000400
#define RIGHT_ALT_PRESSED 0x0001
#define LEFT_ALT_PRESSED 0x0002
#define RIGHT_CTRL_PRESSED 0x0004
#define LEFT_CTRL_PRESSED 0x0008
#define SHIFT_PRESSED 0x0010
#define NUMLOCK_ON 0x0020
#define SCROLLLOCK_ON 0x0040
#define CAPSLOCK_ON 0x0080
#define ENHANCED_KEY 0x0100
#define NLS_DBCSCHAR 0x00010000
#define NLS_ALPHANUMERIC 0x00000000
#define NLS_KATAKANA 0x00020000
#define NLS_HIRAGANA 0x00040000
#define NLS_ROMAN 0x00400000
#define NLS_IME_CONVERSION 0x00800000
#define NLS_IME_DISABLE 0x20000000
#define FROM_LEFT_1ST_BUTTON_PRESSED 0x0001
#define RIGHTMOST_BUTTON_PRESSED 0x0002
#define FROM_LEFT_2ND_BUTTON_PRESSED 0x0004
#define FROM_LEFT_3RD_BUTTON_PRESSED 0x0008
#define FROM_LEFT_4TH_BUTTON_PRESSED 0x0010
#define MOUSE_MOVED 0x0001
#define DOUBLE_CLICK 0x0002
#define MOUSE_WHEELED 0x0004
#define KEY_EVENT 0x0001
#define _MOUSE_EVENT 0x0002
#define WINDOW_BUFFER_SIZE_EVENT 0x0004
#define MENU_EVENT 0x0008
#define FOCUS_EVENT 0x0010
#define FOREGROUND_BLACK 0x0000
#define FOREGROUND_BLUE 0x0001
#define FOREGROUND_GREEN 0x0002
#define FOREGROUND_RED 0x0004
#define FOREGROUND_WHITE 0x0007
#define FOREGROUND_INTENSITY 0x0008
#define BACKGROUND_BLACK 0x0000
#define BACKGROUND_BLUE 0x0010
#define BACKGROUND_GREEN 0x0020
#define BACKGROUND_RED 0x0040
#define BACKGROUND_WHITE 0x0070
#define BACKGROUND_INTENSITY 0x0080
#define COMMON_LVB_LEADING_BYTE 0x0100
#define COMMON_LVB_TRAILING_BYTE 0x0200
#define COMMON_LVB_GRID_HORIZONTAL 0x0400
#define COMMON_LVB_GRID_LVERTICAL 0x0800
#define COMMON_LVB_GRID_RVERTICAL 0x1000
#define COMMON_LVB_REVERSE_VIDEO 0x4000
#define COMMON_LVB_UNDERSCORE 0x8000
#define COMMON_LVB_SBCSDBCS 0x0300
#define CONSOLE_NO_SELECTION 0x0000
#define CONSOLE_SELECTION_IN_PROGRESS 0x0001
#define CONSOLE_SELECTION_NOT_EMPTY 0x0002
#define CONSOLE_MOUSE_SELECTION 0x0004
#define CONSOLE_MOUSE_DOWN 0x0008
#define CTRL_C_EVENT 0
#define CTRL_BREAK_EVENT 1
#define CTRL_CLOSE_EVENT 2
#define CTRL_LOGOFF_EVENT 5
#define CTRL_SHUTDOWN_EVENT 6
#define ENABLE_PROCESSED_INPUT 0x0001
#define ENABLE_LINE_INPUT 0x0002
#define ENABLE_ECHO_INPUT 0x0004
#define ENABLE_WINDOW_INPUT 0x0008
#define ENABLE_MOUSE_INPUT 0x0010
#define ENABLE_PROCESSED_OUTPUT 0x0001
#define ENABLE_WRAP_AT_EOL_OUTPUT 0x0002
#define CONSOLE_TEXTMODE_BUFFER 1
#define MAX_PATH 260
#define HFILE_ERROR -1
#define SYS_WIN32 .T.
#define DLLVER_PLATFORM_NT 0x00000002
#define DLLVER_PLATFORM_WINDOWS 0x00000001
#define FACILITY_WINDOWS 8
#define FACILITY_STORAGE 3
#define FACILITY_RPC 1
#define FACILITY_WIN32 7
#define FACILITY_CONTROL 10
#define FACILITY_NULL 0
#define FACILITY_ITF 4
#define FACILITY_DISPATCH 2
#define ERROR_SUCCESS 0L
#define NO_ERROR 0L
#define ERROR_INVALID_FUNCTION 1L
#define ERROR_FILE_NOT_FOUND 2L
#define ERROR_PATH_NOT_FOUND 3L
#define ERROR_TOO_MANY_OPEN_FILES 4L
#define ERROR_ACCESS_DENIED 5L
#define ERROR_INVALID_HANDLE 6L
#define ERROR_ARENA_TRASHED 7L
#define ERROR_NOT_ENOUGH_MEMORY 8L
#define ERROR_INVALID_BLOCK 9L
#define ERROR_BAD_ENVIRONMENT 10L
#define ERROR_BAD_FORMAT 11L
#define ERROR_INVALID_ACCESS 12L
#define ERROR_INVALID_DATA 13L
#define ERROR_OUTOFMEMORY 14L
#define ERROR_INVALID_DRIVE 15L
#define ERROR_CURRENT_DIRECTORY 16L
#define ERROR_NOT_SAME_DEVICE 17L
#define ERROR_NO_MORE_FILES 18L
#define ERROR_WRITE_PROTECT 19L
#define ERROR_BAD_UNIT 20L
#define ERROR_NOT_READY 21L
#define ERROR_BAD_COMMAND 22L
#define ERROR_CRC 23L
#define ERROR_BAD_LENGTH 24L
#define ERROR_SEEK 25L
#define ERROR_NOT_DOS_DISK 26L
#define ERROR_SECTOR_NOT_FOUND 27L
#define ERROR_OUT_OF_PAPER 28L
#define ERROR_WRITE_FAULT 29L
#define ERROR_READ_FAULT 30L
#define ERROR_GEN_FAILURE 31L
#define ERROR_SHARING_VIOLATION 32L
#define ERROR_LOCK_VIOLATION 33L
#define ERROR_WRONG_DISK 34L
#define ERROR_SHARING_BUFFER_EXCEEDED 36L
#define ERROR_HANDLE_EOF 38L
#define ERROR_HANDLE_DISK_FULL 39L
#define ERROR_NOT_SUPPORTED 50L
#define ERROR_REM_NOT_LIST 51L
#define ERROR_DUP_NAME 52L
#define ERROR_BAD_NETPATH 53L
#define ERROR_NETWORK_BUSY 54L
#define ERROR_DEV_NOT_EXIST 55L
#define ERROR_TOO_MANY_CMDS 56L
#define ERROR_ADAP_HDW_ERR 57L
#define ERROR_BAD_NET_RESP 58L
#define ERROR_UNEXP_NET_ERR 59L
#define ERROR_BAD_REM_ADAP 60L
#define ERROR_PRINTQ_FULL 61L
#define ERROR_NO_SPOOL_SPACE 62L
#define ERROR_PRINT_CANCELLED 63L
#define ERROR_NETNAME_DELETED 64L
#define ERROR_NETWORK_ACCESS_DENIED 65L
#define ERROR_BAD_DEV_TYPE 66L
#define ERROR_BAD_NET_NAME 67L
#define ERROR_TOO_MANY_NAMES 68L
#define ERROR_TOO_MANY_SESS 69L
#define ERROR_SHARING_PAUSED 70L
#define ERROR_REQ_NOT_ACCEP 71L
#define ERROR_REDIR_PAUSED 72L
#define ERROR_FILE_EXISTS 80L
#define ERROR_CANNOT_MAKE 82L
#define ERROR_FAIL_I24 83L
#define ERROR_OUT_OF_STRUCTURES 84L
#define ERROR_ALREADY_ASSIGNED 85L
#define ERROR_INVALID_PASSWORD 86L
#define ERROR_INVALID_PARAMETER 87L
#define ERROR_NET_WRITE_FAULT 88L
#define ERROR_NO_PROC_SLOTS 89L
#define ERROR_TOO_MANY_SEMAPHORES 100L
#define ERROR_EXCL_SEM_ALREADY_OWNED 101L
#define ERROR_SEM_IS_SET 102L
#define ERROR_TOO_MANY_SEM_REQUESTS 103L
#define ERROR_INVALID_AT_INTERRUPT_TIME 104L
#define ERROR_SEM_OWNER_DIED 105L
#define ERROR_SEM_USER_LIMIT 106L
#define ERROR_DISK_CHANGE 107L
#define ERROR_DRIVE_LOCKED 108L
#define ERROR_BROKEN_PIPE 109L
#define ERROR_OPEN_FAILED 110L
#define ERROR_BUFFER_OVERFLOW 111L
#define ERROR_DISK_FULL 112L
#define ERROR_NO_MORE_SEARCH_HANDLES 113L
#define ERROR_INVALID_TARGET_HANDLE 114L
#define ERROR_INVALID_CATEGORY 117L
#define ERROR_INVALID_VERIFY_SWITCH 118L
#define ERROR_BAD_DRIVER_LEVEL 119L
#define ERROR_CALL_NOT_IMPLEMENTED 120L
#define ERROR_SEM_TIMEOUT 121L
#define ERROR_INSUFFICIENT_BUFFER 122L
#define ERROR_INVALID_NAME 123L
#define ERROR_INVALID_LEVEL 124L
#define ERROR_NO_VOLUME_LABEL 125L
#define ERROR_MOD_NOT_FOUND 126L
#define ERROR_PROC_NOT_FOUND 127L
#define ERROR_WAIT_NO_CHILDREN 128L
#define ERROR_CHILD_NOT_COMPLETE 129L
#define ERROR_DIRECT_ACCESS_HANDLE 130L
#define ERROR_NEGATIVE_SEEK 131L
#define ERROR_SEEK_ON_DEVICE 132L
#define ERROR_IS_JOIN_TARGET 133L
#define ERROR_IS_JOINED 134L
#define ERROR_IS_SUBSTED 135L
#define ERROR_NOT_JOINED 136L
#define ERROR_NOT_SUBSTED 137L
#define ERROR_JOIN_TO_JOIN 138L
#define ERROR_SUBST_TO_SUBST 139L
#define ERROR_JOIN_TO_SUBST 140L
#define ERROR_SUBST_TO_JOIN 141L
#define ERROR_BUSY_DRIVE 142L
#define ERROR_SAME_DRIVE 143L
#define ERROR_DIR_NOT_ROOT 144L
#define ERROR_DIR_NOT_EMPTY 145L
#define ERROR_IS_SUBST_PATH 146L
#define ERROR_IS_JOIN_PATH 147L
#define ERROR_PATH_BUSY 148L
#define ERROR_IS_SUBST_TARGET 149L
#define ERROR_SYSTEM_TRACE 150L
#define ERROR_INVALID_EVENT_COUNT 151L
#define ERROR_TOO_MANY_MUXWAITERS 152L
#define ERROR_INVALID_LIST_FORMAT 153L
#define ERROR_LABEL_TOO_LONG 154L
#define ERROR_TOO_MANY_TCBS 155L
#define ERROR_SIGNAL_REFUSED 156L
#define ERROR_DISCARDED 157L
#define ERROR_NOT_LOCKED 158L
#define ERROR_BAD_THREADID_ADDR 159L
#define ERROR_BAD_ARGUMENTS 160L
#define ERROR_BAD_PATHNAME 161L
#define ERROR_SIGNAL_PENDING 162L
#define ERROR_MAX_THRDS_REACHED 164L
#define ERROR_LOCK_FAILED 167L
#define ERROR_BUSY 170L
#define ERROR_CANCEL_VIOLATION 173L
#define ERROR_ATOMIC_LOCKS_NOT_SUPPORTED 174L
#define ERROR_INVALID_SEGMENT_NUMBER 180L
#define ERROR_INVALID_ORDINAL 182L
#define ERROR_ALREADY_EXISTS 183L
#define ERROR_INVALID_FLAG_NUMBER 186L
#define ERROR_SEM_NOT_FOUND 187L
#define ERROR_INVALID_STARTING_CODESEG 188L
#define ERROR_INVALID_STACKSEG 189L
#define ERROR_INVALID_MODULETYPE 190L
#define ERROR_INVALID_EXE_SIGNATURE 191L
#define ERROR_EXE_MARKED_INVALID 192L
#define ERROR_BAD_EXE_FORMAT 193L
#define ERROR_ITERATED_DATA_EXCEEDS_64k 194L
#define ERROR_INVALID_MINALLOCSIZE 195L
#define ERROR_DYNLINK_FROM_INVALID_RING 196L
#define ERROR_IOPL_NOT_ENABLED 197L
#define ERROR_INVALID_SEGDPL 198L
#define ERROR_AUTODATASEG_EXCEEDS_64k 199L
#define ERROR_RING2SEG_MUST_BE_MOVABLE 200L
#define ERROR_RELOC_CHAIN_XEEDS_SEGLIM 201L
#define ERROR_INFLOOP_IN_RELOC_CHAIN 202L
#define ERROR_ENVVAR_NOT_FOUND 203L
#define ERROR_NO_SIGNAL_SENT 205L
#define ERROR_FILENAME_EXCED_RANGE 206L
#define ERROR_RING2_STACK_IN_USE 207L
#define ERROR_META_EXPANSION_TOO_LONG 208L
#define ERROR_INVALID_SIGNAL_NUMBER 209L
#define ERROR_THREAD_1_INACTIVE 210L
#define ERROR_LOCKED 212L
#define ERROR_TOO_MANY_MODULES 214L
#define ERROR_NESTING_NOT_ALLOWED 215L
#define ERROR_BAD_PIPE 230L
#define ERROR_PIPE_BUSY 231L
#define ERROR_NO_DATA 232L
#define ERROR_PIPE_NOT_CONNECTED 233L
#define ERROR_MORE_DATA 234L
#define ERROR_VC_DISCONNECTED 240L
#define ERROR_INVALID_EA_NAME 254L
#define ERROR_EA_LIST_INCONSISTENT 255L
#define ERROR_NO_MORE_ITEMS 259L
#define ERROR_CANNOT_COPY 266L
#define ERROR_DIRECTORY 267L
#define ERROR_EAS_DIDNT_FIT 275L
#define ERROR_EA_FILE_CORRUPT 276L
#define ERROR_EA_TABLE_FULL 277L
#define ERROR_INVALID_EA_HANDLE 278L
#define ERROR_EAS_NOT_SUPPORTED 282L
#define ERROR_NOT_OWNER 288L
#define ERROR_TOO_MANY_POSTS 298L
#define ERROR_PARTIAL_COPY 299L
#define ERROR_MR_MID_NOT_FOUND 317L
#define ERROR_INVALID_ADDRESS 487L
#define ERROR_ARITHMETIC_OVERFLOW 534L
#define ERROR_PIPE_CONNECTED 535L
#define ERROR_PIPE_LISTENING 536L
#define ERROR_EA_ACCESS_DENIED 994L
#define ERROR_OPERATION_ABORTED 995L
#define ERROR_IO_INCOMPLETE 996L
#define ERROR_IO_PENDING 997L
#define ERROR_NOACCESS 998L
#define ERROR_SWAPERROR 999L
#define ERROR_STACK_OVERFLOW 1001L
#define ERROR_INVALID_MESSAGE 1002L
#define ERROR_CAN_NOT_COMPLETE 1003L
#define ERROR_INVALID_FLAGS 1004L
#define ERROR_UNRECOGNIZED_VOLUME 1005L
#define ERROR_FILE_INVALID 1006L
#define ERROR_FULLSCREEN_MODE 1007L
#define ERROR_NO_TOKEN 1008L
#define ERROR_BADDB 1009L
#define ERROR_BADKEY 1010L
#define ERROR_CANTOPEN 1011L
#define ERROR_CANTREAD 1012L
#define ERROR_CANTWRITE 1013L
#define ERROR_REGISTRY_RECOVERED 1014L
#define ERROR_REGISTRY_CORRUPT 1015L
#define ERROR_REGISTRY_IO_FAILED 1016L
#define ERROR_NOT_REGISTRY_FILE 1017L
#define ERROR_KEY_DELETED 1018L
#define ERROR_NO_LOG_SPACE 1019L
#define ERROR_KEY_HAS_CHILDREN 1020L
#define ERROR_CHILD_MUST_BE_VOLATILE 1021L
#define ERROR_NOTIFY_ENUM_DIR 1022L
#define ERROR_DEPENDENT_SERVICES_RUNNING 1051L
#define ERROR_INVALID_SERVICE_CONTROL 1052L
#define ERROR_SERVICE_REQUEST_TIMEOUT 1053L
#define ERROR_SERVICE_NO_THREAD 1054L
#define ERROR_SERVICE_DATABASE_LOCKED 1055L
#define ERROR_SERVICE_ALREADY_RUNNING 1056L
#define ERROR_INVALID_SERVICE_ACCOUNT 1057L
#define ERROR_SERVICE_DISABLED 1058L
#define ERROR_CIRCULAR_DEPENDENCY 1059L
#define ERROR_SERVICE_DOES_NOT_EXIST 1060L
#define ERROR_SERVICE_CANNOT_ACCEPT_CTRL 1061L
#define ERROR_SERVICE_NOT_ACTIVE 1062L
#define ERROR_FAILED_SERVICE_CONTROLLER_CONNECT 1063L
#define ERROR_EXCEPTION_IN_SERVICE 1064L
#define ERROR_DATABASE_DOES_NOT_EXIST 1065L
#define ERROR_SERVICE_SPECIFIC_ERROR 1066L
#define ERROR_PROCESS_ABORTED 1067L
#define ERROR_SERVICE_DEPENDENCY_FAIL 1068L
#define ERROR_SERVICE_LOGON_FAILED 1069L
#define ERROR_SERVICE_START_HANG 1070L
#define ERROR_INVALID_SERVICE_LOCK 1071L
#define ERROR_SERVICE_MARKED_FOR_DELETE 1072L
#define ERROR_SERVICE_EXISTS 1073L
#define ERROR_ALREADY_RUNNING_LKG 1074L
#define ERROR_SERVICE_DEPENDENCY_DELETED 1075L
#define ERROR_BOOT_ALREADY_ACCEPTED 1076L
#define ERROR_SERVICE_NEVER_STARTED 1077L
#define ERROR_DUPLICATE_SERVICE_NAME 1078L
#define ERROR_END_OF_MEDIA 1100L
#define ERROR_FILEMARK_DETECTED 1101L
#define ERROR_BEGINNING_OF_MEDIA 1102L
#define ERROR_SETMARK_DETECTED 1103L
#define ERROR_NO_DATA_DETECTED 1104L
#define ERROR_PARTITION_FAILURE 1105L
#define ERROR_INVALID_BLOCK_LENGTH 1106L
#define ERROR_DEVICE_NOT_PARTITIONED 1107L
#define ERROR_UNABLE_TO_LOCK_MEDIA 1108L
#define ERROR_UNABLE_TO_UNLOAD_MEDIA 1109L
#define ERROR_MEDIA_CHANGED 1110L
#define ERROR_BUS_RESET 1111L
#define ERROR_NO_MEDIA_IN_DRIVE 1112L
#define ERROR_NO_UNICODE_TRANSLATION 1113L
#define ERROR_DLL_INIT_FAILED 1114L
#define ERROR_SHUTDOWN_IN_PROGRESS 1115L
#define ERROR_NO_SHUTDOWN_IN_PROGRESS 1116L
#define ERROR_IO_DEVICE 1117L
#define ERROR_SERIAL_NO_DEVICE 1118L
#define ERROR_IRQ_BUSY 1119L
#define ERROR_MORE_WRITES 1120L
#define ERROR_COUNTER_TIMEOUT 1121L
#define ERROR_FLOPPY_ID_MARK_NOT_FOUND 1122L
#define ERROR_FLOPPY_WRONG_CYLINDER 1123L
#define ERROR_FLOPPY_UNKNOWN_ERROR 1124L
#define ERROR_FLOPPY_BAD_REGISTERS 1125L
#define ERROR_DISK_RECALIBRATE_FAILED 1126L
#define ERROR_DISK_OPERATION_FAILED 1127L
#define ERROR_DISK_RESET_FAILED 1128L
#define ERROR_EOM_OVERFLOW 1129L
#define ERROR_NOT_ENOUGH_SERVER_MEMORY 1130L
#define ERROR_POSSIBLE_DEADLOCK 1131L
#define ERROR_MAPPED_ALIGNMENT 1132L
#define ERROR_SET_POWER_STATE_VETOED 1140L
#define ERROR_SET_POWER_STATE_FAILED 1141L
#define ERROR_OLD_WIN_VERSION 1150L
#define ERROR_APP_WRONG_OS 1151L
#define ERROR_SINGLE_INSTANCE_APP 1152L
#define ERROR_RMODE_APP 1153L
#define ERROR_INVALID_DLL 1154L
#define ERROR_NO_ASSOCIATION 1155L
#define ERROR_DDE_FAIL 1156L
#define ERROR_DLL_NOT_FOUND 1157L
#define ERROR_BAD_USERNAME 2202L
#define ERROR_NOT_CONNECTED 2250L
#define ERROR_OPEN_FILES 2401L
#define ERROR_ACTIVE_CONNECTIONS 2402L
#define ERROR_DEVICE_IN_USE 2404L
#define ERROR_BAD_DEVICE 1200L
#define ERROR_CONNECTION_UNAVAIL 1201L
#define ERROR_DEVICE_ALREADY_REMEMBERED 1202L
#define ERROR_NO_NET_OR_BAD_PATH 1203L
#define ERROR_BAD_PROVIDER 1204L
#define ERROR_CANNOT_OPEN_PROFILE 1205L
#define ERROR_BAD_PROFILE 1206L
#define ERROR_NOT_CONTAINER 1207L
#define ERROR_EXTENDED_ERROR 1208L
#define ERROR_INVALID_GROUPNAME 1209L
#define ERROR_INVALID_COMPUTERNAME 1210L
#define ERROR_INVALID_EVENTNAME 1211L
#define ERROR_INVALID_DOMAINNAME 1212L
#define ERROR_INVALID_SERVICENAME 1213L
#define ERROR_INVALID_NETNAME 1214L
#define ERROR_INVALID_SHARENAME 1215L
#define ERROR_INVALID_PASSWORDNAME 1216L
#define ERROR_INVALID_MESSAGENAME 1217L
#define ERROR_INVALID_MESSAGEDEST 1218L
#define ERROR_SESSION_CREDENTIAL_CONFLICT 1219L
#define ERROR_REMOTE_SESSION_LIMIT_EXCEEDED 1220L
#define ERROR_DUP_DOMAINNAME 1221L
#define ERROR_NO_NETWORK 1222L
#define ERROR_CANCELLED 1223L
#define ERROR_USER_MAPPED_FILE 1224L
#define ERROR_CONNECTION_REFUSED 1225L
#define ERROR_GRACEFUL_DISCONNECT 1226L
#define ERROR_ADDRESS_ALREADY_ASSOCIATED 1227L
#define ERROR_ADDRESS_NOT_ASSOCIATED 1228L
#define ERROR_CONNECTION_INVALID 1229L
#define ERROR_CONNECTION_ACTIVE 1230L
#define ERROR_NETWORK_UNREACHABLE 1231L
#define ERROR_HOST_UNREACHABLE 1232L
#define ERROR_PROTOCOL_UNREACHABLE 1233L
#define ERROR_PORT_UNREACHABLE 1234L
#define ERROR_REQUEST_ABORTED 1235L
#define ERROR_CONNECTION_ABORTED 1236L
#define ERROR_RETRY 1237L
#define ERROR_CONNECTION_COUNT_LIMIT 1238L
#define ERROR_LOGIN_TIME_RESTRICTION 1239L
#define ERROR_LOGIN_WKSTA_RESTRICTION 1240L
#define ERROR_INCORRECT_ADDRESS 1241L
#define ERROR_ALREADY_REGISTERED 1242L
#define ERROR_SERVICE_NOT_FOUND 1243L
#define ERROR_NOT_AUTHENTICATED 1244L
#define ERROR_NOT_LOGGED_ON 1245L
#define ERROR_CONTINUE 1246L
#define ERROR_ALREADY_INITIALIZED 1247L
#define ERROR_NO_MORE_DEVICES 1248L
#define ERROR_NOT_ALL_ASSIGNED 1300L
#define ERROR_SOME_NOT_MAPPED 1301L
#define ERROR_NO_QUOTAS_FOR_ACCOUNT 1302L
#define ERROR_LOCAL_USER_SESSION_KEY 1303L
#define ERROR_NULL_LM_PASSWORD 1304L
#define ERROR_UNKNOWN_REVISION 1305L
#define ERROR_REVISION_MISMATCH 1306L
#define ERROR_INVALID_OWNER 1307L
#define ERROR_INVALID_PRIMARY_GROUP 1308L
#define ERROR_NO_IMPERSONATION_TOKEN 1309L
#define ERROR_CANT_DISABLE_MANDATORY 1310L
#define ERROR_NO_LOGON_SERVERS 1311L
#define ERROR_NO_SUCH_LOGON_SESSION 1312L
#define ERROR_NO_SUCH_PRIVILEGE 1313L
#define ERROR_PRIVILEGE_NOT_HELD 1314L
#define ERROR_INVALID_ACCOUNT_NAME 1315L
#define ERROR_USER_EXISTS 1316L
#define ERROR_NO_SUCH_USER 1317L
#define ERROR_GROUP_EXISTS 1318L
#define ERROR_NO_SUCH_GROUP 1319L
#define ERROR_MEMBER_IN_GROUP 1320L
#define ERROR_MEMBER_NOT_IN_GROUP 1321L
#define ERROR_LAST_ADMIN 1322L
#define ERROR_WRONG_PASSWORD 1323L
#define ERROR_ILL_FORMED_PASSWORD 1324L
#define ERROR_PASSWORD_RESTRICTION 1325L
#define ERROR_LOGON_FAILURE 1326L
#define ERROR_ACCOUNT_RESTRICTION 1327L
#define ERROR_INVALID_LOGON_HOURS 1328L
#define ERROR_INVALID_WORKSTATION 1329L
#define ERROR_PASSWORD_EXPIRED 1330L
#define ERROR_ACCOUNT_DISABLED 1331L
#define ERROR_NONE_MAPPED 1332L
#define ERROR_TOO_MANY_LUIDS_REQUESTED 1333L
#define ERROR_LUIDS_EXHAUSTED 1334L
#define ERROR_INVALID_SUB_AUTHORITY 1335L
#define ERROR_INVALID_ACL 1336L
#define ERROR_INVALID_SID 1337L
#define ERROR_INVALID_SECURITY_DESCR 1338L
#define ERROR_BAD_INHERITANCE_ACL 1340L
#define ERROR_SERVER_DISABLED 1341L
#define ERROR_SERVER_NOT_DISABLED 1342L
#define ERROR_INVALID_ID_AUTHORITY 1343L
#define ERROR_ALLOTTED_SPACE_EXCEEDED 1344L
#define ERROR_INVALID_GROUP_ATTRIBUTES 1345L
#define ERROR_BAD_IMPERSONATION_LEVEL 1346L
#define ERROR_CANT_OPEN_ANONYMOUS 1347L
#define ERROR_BAD_VALIDATION_CLASS 1348L
#define ERROR_BAD_TOKEN_TYPE 1349L
#define ERROR_NO_SECURITY_ON_OBJECT 1350L
#define ERROR_CANT_ACCESS_DOMAIN_INFO 1351L
#define ERROR_INVALID_SERVER_STATE 1352L
#define ERROR_INVALID_DOMAIN_STATE 1353L
#define ERROR_INVALID_DOMAIN_ROLE 1354L
#define ERROR_NO_SUCH_DOMAIN 1355L
#define ERROR_DOMAIN_EXISTS 1356L
#define ERROR_DOMAIN_LIMIT_EXCEEDED 1357L
#define ERROR_INTERNAL_DB_CORRUPTION 1358L
#define ERROR_INTERNAL_ERROR 1359L
#define ERROR_GENERIC_NOT_MAPPED 1360L
#define ERROR_BAD_DESCRIPTOR_FORMAT 1361L
#define ERROR_NOT_LOGON_PROCESS 1362L
#define ERROR_LOGON_SESSION_EXISTS 1363L
#define ERROR_NO_SUCH_PACKAGE 1364L
#define ERROR_BAD_LOGON_SESSION_STATE 1365L
#define ERROR_LOGON_SESSION_COLLISION 1366L
#define ERROR_INVALID_LOGON_TYPE 1367L
#define ERROR_CANNOT_IMPERSONATE 1368L
#define ERROR_RXACT_INVALID_STATE 1369L
#define ERROR_RXACT_COMMIT_FAILURE 1370L
#define ERROR_SPECIAL_ACCOUNT 1371L
#define ERROR_SPECIAL_GROUP 1372L
#define ERROR_SPECIAL_USER 1373L
#define ERROR_MEMBERS_PRIMARY_GROUP 1374L
#define ERROR_TOKEN_ALREADY_IN_USE 1375L
#define ERROR_NO_SUCH_ALIAS 1376L
#define ERROR_MEMBER_NOT_IN_ALIAS 1377L
#define ERROR_MEMBER_IN_ALIAS 1378L
#define ERROR_ALIAS_EXISTS 1379L
#define ERROR_LOGON_NOT_GRANTED 1380L
#define ERROR_TOO_MANY_SECRETS 1381L
#define ERROR_SECRET_TOO_LONG 1382L
#define ERROR_INTERNAL_DB_ERROR 1383L
#define ERROR_TOO_MANY_CONTEXT_IDS 1384L
#define ERROR_LOGON_TYPE_NOT_GRANTED 1385L
#define ERROR_NT_CROSS_ENCRYPTION_REQUIRED 1386L
#define ERROR_NO_SUCH_MEMBER 1387L
#define ERROR_INVALID_MEMBER 1388L
#define ERROR_TOO_MANY_SIDS 1389L
#define ERROR_LM_CROSS_ENCRYPTION_REQUIRED 1390L
#define ERROR_NO_INHERITANCE 1391L
#define ERROR_FILE_CORRUPT 1392L
#define ERROR_DISK_CORRUPT 1393L
#define ERROR_NO_USER_SESSION_KEY 1394L
#define ERROR_LICENSE_QUOTA_EXCEEDED 1395L
#define ERROR_INVALID_WINDOW_HANDLE 1400L
#define ERROR_INVALID_MENU_HANDLE 1401L
#define ERROR_INVALID_CURSOR_HANDLE 1402L
#define ERROR_INVALID_ACCEL_HANDLE 1403L
#define ERROR_INVALID_HOOK_HANDLE 1404L
#define ERROR_INVALID_DWP_HANDLE 1405L
#define ERROR_TLW_WITH_WSCHILD 1406L
#define ERROR_CANNOT_FIND_WND_CLASS 1407L
#define ERROR_WINDOW_OF_OTHER_THREAD 1408L
#define ERROR_HOTKEY_ALREADY_REGISTERED 1409L
#define ERROR_CLASS_ALREADY_EXISTS 1410L
#define ERROR_CLASS_DOES_NOT_EXIST 1411L
#define ERROR_CLASS_HAS_WINDOWS 1412L
#define ERROR_INVALID_INDEX 1413L
#define ERROR_INVALID_ICON_HANDLE 1414L
#define ERROR_PRIVATE_DIALOG_INDEX 1415L
#define ERROR_LISTBOX_ID_NOT_FOUND 1416L
#define ERROR_NO_WILDCARD_CHARACTERS 1417L
#define ERROR_CLIPBOARD_NOT_OPEN 1418L
#define ERROR_HOTKEY_NOT_REGISTERED 1419L
#define ERROR_WINDOW_NOT_DIALOG 1420L
#define ERROR_CONTROL_ID_NOT_FOUND 1421L
#define ERROR_INVALID_COMBOBOX_MESSAGE 1422L
#define ERROR_WINDOW_NOT_COMBOBOX 1423L
#define ERROR_INVALID_EDIT_HEIGHT 1424L
#define ERROR_DC_NOT_FOUND 1425L
#define ERROR_INVALID_HOOK_FILTER 1426L
#define ERROR_INVALID_FILTER_PROC 1427L
#define ERROR_HOOK_NEEDS_HMOD 1428L
#define ERROR_GLOBAL_ONLY_HOOK 1429L
#define ERROR_JOURNAL_HOOK_SET 1430L
#define ERROR_HOOK_NOT_INSTALLED 1431L
#define ERROR_INVALID_LB_MESSAGE 1432L
#define ERROR_SETCOUNT_ON_BAD_LB 1433L
#define ERROR_LB_WITHOUT_TABSTOPS 1434L
#define ERROR_DESTROY_OBJECT_OF_OTHER_THREAD 1435L
#define ERROR_CHILD_WINDOW_MENU 1436L
#define ERROR_NO_SYSTEM_MENU 1437L
#define ERROR_INVALID_MSGBOX_STYLE 1438L
#define ERROR_INVALID_SPI_VALUE 1439L
#define ERROR_SCREEN_ALREADY_LOCKED 1440L
#define ERROR_HWNDS_HAVE_DIFF_PARENT 1441L
#define ERROR_NOT_CHILD_WINDOW 1442L
#define ERROR_INVALID_GW_COMMAND 1443L
#define ERROR_INVALID_THREAD_ID 1444L
#define ERROR_NON_MDICHILD_WINDOW 1445L
#define ERROR_POPUP_ALREADY_ACTIVE 1446L
#define ERROR_NO_SCROLLBARS 1447L
#define ERROR_INVALID_SCROLLBAR_RANGE 1448L
#define ERROR_INVALID_SHOWWIN_COMMAND 1449L
#define ERROR_NO_SYSTEM_RESOURCES 1450L
#define ERROR_NONPAGED_SYSTEM_RESOURCES 1451L
#define ERROR_PAGED_SYSTEM_RESOURCES 1452L
#define ERROR_WORKING_SET_QUOTA 1453L
#define ERROR_PAGEFILE_QUOTA 1454L
#define ERROR_COMMITMENT_LIMIT 1455L
#define ERROR_MENU_ITEM_NOT_FOUND 1456L
#define ERROR_EVENTLOG_FILE_CORRUPT 1500L
#define ERROR_EVENTLOG_CANT_START 1501L
#define ERROR_LOG_FILE_FULL 1502L
#define ERROR_EVENTLOG_FILE_CHANGED 1503L
#define RPC_S_INVALID_STRING_BINDING 1700L
#define RPC_S_WRONG_KIND_OF_BINDING 1701L
#define RPC_S_INVALID_BINDING 1702L
#define RPC_S_PROTSEQ_NOT_SUPPORTED 1703L
#define RPC_S_INVALID_RPC_PROTSEQ 1704L
#define RPC_S_INVALID_STRING_UUID 1705L
#define RPC_S_INVALID_ENDPOINT_FORMAT 1706L
#define RPC_S_INVALID_NET_ADDR 1707L
#define RPC_S_NO_ENDPOINT_FOUND 1708L
#define RPC_S_INVALID_TIMEOUT 1709L
#define RPC_S_OBJECT_NOT_FOUND 1710L
#define RPC_S_ALREADY_REGISTERED 1711L
#define RPC_S_TYPE_ALREADY_REGISTERED 1712L
#define RPC_S_ALREADY_LISTENING 1713L
#define RPC_S_NO_PROTSEQS_REGISTERED 1714L
#define RPC_S_NOT_LISTENING 1715L
#define RPC_S_UNKNOWN_MGR_TYPE 1716L
#define RPC_S_UNKNOWN_IF 1717L
#define RPC_S_NO_BINDINGS 1718L
#define RPC_S_NO_PROTSEQS 1719L
#define RPC_S_CANT_CREATE_ENDPOINT 1720L
#define RPC_S_OUT_OF_RESOURCES 1721L
#define RPC_S_SERVER_UNAVAILABLE 1722L
#define RPC_S_SERVER_TOO_BUSY 1723L
#define RPC_S_INVALID_NETWORK_OPTIONS 1724L
#define RPC_S_NO_CALL_ACTIVE 1725L
#define RPC_S_CALL_FAILED 1726L
#define RPC_S_CALL_FAILED_DNE 1727L
#define RPC_S_PROTOCOL_ERROR 1728L
#define RPC_S_UNSUPPORTED_TRANS_SYN 1730L
#define RPC_S_UNSUPPORTED_TYPE 1732L
#define RPC_S_INVALID_TAG 1733L
#define RPC_S_INVALID_BOUND 1734L
#define RPC_S_NO_ENTRY_NAME 1735L
#define RPC_S_INVALID_NAME_SYNTAX 1736L
#define RPC_S_UNSUPPORTED_NAME_SYNTAX 1737L
#define RPC_S_UUID_NO_ADDRESS 1739L
#define RPC_S_DUPLICATE_ENDPOINT 1740L
#define RPC_S_UNKNOWN_AUTHN_TYPE 1741L
#define RPC_S_MAX_CALLS_TOO_SMALL 1742L
#define RPC_S_STRING_TOO_LONG 1743L
#define RPC_S_PROTSEQ_NOT_FOUND 1744L
#define RPC_S_PROCNUM_OUT_OF_RANGE 1745L
#define RPC_S_BINDING_HAS_NO_AUTH 1746L
#define RPC_S_UNKNOWN_AUTHN_SERVICE 1747L
#define RPC_S_UNKNOWN_AUTHN_LEVEL 1748L
#define RPC_S_INVALID_AUTH_IDENTITY 1749L
#define RPC_S_UNKNOWN_AUTHZ_SERVICE 1750L
#define EPT_S_INVALID_ENTRY 1751L
#define EPT_S_CANT_PERFORM_OP 1752L
#define EPT_S_NOT_REGISTERED 1753L
#define RPC_S_NOTHING_TO_EXPORT 1754L
#define RPC_S_INCOMPLETE_NAME 1755L
#define RPC_S_INVALID_VERS_OPTION 1756L
#define RPC_S_NO_MORE_MEMBERS 1757L
#define RPC_S_NOT_ALL_OBJS_UNEXPORTED 1758L
#define RPC_S_INTERFACE_NOT_FOUND 1759L
#define RPC_S_ENTRY_ALREADY_EXISTS 1760L
#define RPC_S_ENTRY_NOT_FOUND 1761L
#define RPC_S_NAME_SERVICE_UNAVAILABLE 1762L
#define RPC_S_INVALID_NAF_ID 1763L
#define RPC_S_CANNOT_SUPPORT 1764L
#define RPC_S_NO_CONTEXT_AVAILABLE 1765L
#define RPC_S_INTERNAL_ERROR 1766L
#define RPC_S_ZERO_DIVIDE 1767L
#define RPC_S_ADDRESS_ERROR 1768L
#define RPC_S_FP_DIV_ZERO 1769L
#define RPC_S_FP_UNDERFLOW 1770L
#define RPC_S_FP_OVERFLOW 1771L
#define RPC_X_NO_MORE_ENTRIES 1772L
#define RPC_X_SS_CHAR_TRANS_OPEN_FAIL 1773L
#define RPC_X_SS_CHAR_TRANS_SHORT_FILE 1774L
#define RPC_X_SS_IN_NULL_CONTEXT 1775L
#define RPC_X_SS_CONTEXT_DAMAGED 1777L
#define RPC_X_SS_HANDLES_MISMATCH 1778L
#define RPC_X_SS_CANNOT_GET_CALL_HANDLE 1779L
#define RPC_X_NULL_REF_POINTER 1780L
#define RPC_X_ENUM_VALUE_OUT_OF_RANGE 1781L
#define RPC_X_BYTE_COUNT_TOO_SMALL 1782L
#define RPC_X_BAD_STUB_DATA 1783L
#define ERROR_INVALID_USER_BUFFER 1784L
#define ERROR_UNRECOGNIZED_MEDIA 1785L
#define ERROR_NO_TRUST_LSA_SECRET 1786L
#define ERROR_NO_TRUST_SAM_ACCOUNT 1787L
#define ERROR_TRUSTED_DOMAIN_FAILURE 1788L
#define ERROR_TRUSTED_RELATIONSHIP_FAILURE 1789L
#define ERROR_TRUST_FAILURE 1790L
#define RPC_S_CALL_IN_PROGRESS 1791L
#define ERROR_NETLOGON_NOT_STARTED 1792L
#define ERROR_ACCOUNT_EXPIRED 1793L
#define ERROR_REDIRECTOR_HAS_OPEN_HANDLES 1794L
#define ERROR_PRINTER_DRIVER_ALREADY_INSTALLED 1795L
#define ERROR_UNKNOWN_PORT 1796L
#define ERROR_UNKNOWN_PRINTER_DRIVER 1797L
#define ERROR_UNKNOWN_PRINTPROCESSOR 1798L
#define ERROR_INVALID_SEPARATOR_FILE 1799L
#define ERROR_INVALID_PRIORITY 1800L
#define ERROR_INVALID_PRINTER_NAME 1801L
#define ERROR_PRINTER_ALREADY_EXISTS 1802L
#define ERROR_INVALID_PRINTER_COMMAND 1803L
#define ERROR_INVALID_DATATYPE 1804L
#define ERROR_INVALID_ENVIRONMENT 1805L
#define RPC_S_NO_MORE_BINDINGS 1806L
#define ERROR_NOLOGON_INTERDOMAIN_TRUST_ACCOUNT 1807L
#define ERROR_NOLOGON_WORKSTATION_TRUST_ACCOUNT 1808L
#define ERROR_NOLOGON_SERVER_TRUST_ACCOUNT 1809L
#define ERROR_DOMAIN_TRUST_INCONSISTENT 1810L
#define ERROR_SERVER_HAS_OPEN_HANDLES 1811L
#define ERROR_RESOURCE_DATA_NOT_FOUND 1812L
#define ERROR_RESOURCE_TYPE_NOT_FOUND 1813L
#define ERROR_RESOURCE_NAME_NOT_FOUND 1814L
#define ERROR_RESOURCE_LANG_NOT_FOUND 1815L
#define ERROR_NOT_ENOUGH_QUOTA 1816L
#define RPC_S_NO_INTERFACES 1817L
#define RPC_S_CALL_CANCELLED 1818L
#define RPC_S_BINDING_INCOMPLETE 1819L
#define RPC_S_COMM_FAILURE 1820L
#define RPC_S_UNSUPPORTED_AUTHN_LEVEL 1821L
#define RPC_S_NO_PRINC_NAME 1822L
#define RPC_S_NOT_RPC_ERROR 1823L
#define RPC_S_UUID_LOCAL_ONLY 1824L
#define RPC_S_SEC_PKG_ERROR 1825L
#define RPC_S_NOT_CANCELLED 1826L
#define RPC_X_INVALID_ES_ACTION 1827L
#define RPC_X_WRONG_ES_VERSION 1828L
#define RPC_X_WRONG_STUB_VERSION 1829L
#define RPC_S_GROUP_MEMBER_NOT_FOUND 1898L
#define EPT_S_CANT_CREATE 1899L
#define RPC_S_INVALID_OBJECT 1900L
#define ERROR_INVALID_TIME 1901L
#define ERROR_INVALID_FORM_NAME 1902L
#define ERROR_INVALID_FORM_SIZE 1903L
#define ERROR_ALREADY_WAITING 1904L
#define ERROR_PRINTER_DELETED 1905L
#define ERROR_INVALID_PRINTER_STATE 1906L
#define ERROR_PASSWORD_MUST_CHANGE 1907L
#define ERROR_DOMAIN_CONTROLLER_NOT_FOUND 1908L
#define ERROR_ACCOUNT_LOCKED_OUT 1909L
#define ERROR_NO_BROWSER_SERVERS_FOUND 6118L
#define ERROR_INVALID_PIXEL_FORMAT 2000L
#define ERROR_BAD_DRIVER 2001L
#define ERROR_INVALID_WINDOW_STYLE 2002L
#define ERROR_METAFILE_NOT_SUPPORTED 2003L
#define ERROR_TRANSFORM_NOT_SUPPORTED 2004L
#define ERROR_CLIPPING_NOT_SUPPORTED 2005L
#define ERROR_UNKNOWN_PRINT_MONITOR 3000L
#define ERROR_PRINTER_DRIVER_IN_USE 3001L
#define ERROR_SPOOL_FILE_NOT_FOUND 3002L
#define ERROR_SPL_NO_STARTDOC 3003L
#define ERROR_SPL_NO_ADDJOB 3004L
#define ERROR_PRINT_PROCESSOR_ALREADY_INSTALLED 3005L
#define ERROR_PRINT_MONITOR_ALREADY_INSTALLED 3006L
#define ERROR_WINS_INTERNAL 4000L
#define ERROR_CAN_NOT_DEL_LOCAL_WINS 4001L
#define ERROR_STATIC_INIT 4002L
#define ERROR_INC_BACKUP 4003L
#define ERROR_FULL_BACKUP 4004L
#define ERROR_REC_NON_EXISTENT 4005L
#define ERROR_RPL_NOT_ALLOWED 4006L
#define SEVERITY_SUCCESS 0
#define SEVERITY_ERROR 1
#define FACILITY_NT_BIT 0x10000000
#define S_OK 0x00000000L
#define NOERROR S_OK
#define E_UNEXPECTED 0x8000FFFFL
#define E_NOTIMPL 0x80004001L
#define E_OUTOFMEMORY 0x8007000EL
#define E_INVALIDARG 0x80070057L
#define E_NOINTERFACE 0x80004002L
#define E_POINTER 0x80004003L
#define E_HANDLE 0x80070006L
#define E_ABORT 0x80004004L
#define E_FAIL 0x80004005L
#define E_ACCESSDENIED 0x80070005L
#define CO_E_INIT_TLS 0x80004006L
#define CO_E_INIT_SHARED_ALLOCATOR 0x80004007L
#define CO_E_INIT_MEMORY_ALLOCATOR 0x80004008L
#define CO_E_INIT_CLASS_CACHE 0x80004009L
#define CO_E_INIT_RPC_CHANNEL 0x8000400AL
#define CO_E_INIT_TLS_SET_CHANNEL_CONTROL 0x8000400BL
#define CO_E_INIT_TLS_CHANNEL_CONTROL 0x8000400CL
#define CO_E_INIT_UNACCEPTED_USER_ALLOCATOR 0x8000400DL
#define CO_E_INIT_SCM_MUTEX_EXISTS 0x8000400EL
#define CO_E_INIT_SCM_FILE_MAPPING_EXISTS 0x8000400FL
#define CO_E_INIT_SCM_MAP_VIEW_OF_FILE 0x80004010L
#define CO_E_INIT_SCM_EXEC_FAILURE 0x80004011L
#define CO_E_INIT_ONLY_SINGLE_THREADED 0x80004012L
#define S_FALSE 0x00000001L
#define OLE_E_FIRST 0x80040000L
#define OLE_E_LAST 0x800400FFL
#define OLE_S_FIRST 0x00040000L
#define OLE_S_LAST 0x000400FFL
#define OLE_E_OLEVERB 0x80040000L
#define OLE_E_ADVF 0x80040001L
#define OLE_E_ENUM_NOMORE 0x80040002L
#define OLE_E_ADVISENOTSUPPORTED 0x80040003L
#define OLE_E_NOCONNECTION 0x80040004L
#define OLE_E_NOTRUNNING 0x80040005L
#define OLE_E_NOCACHE 0x80040006L
#define OLE_E_BLANK 0x80040007L
#define OLE_E_CLASSDIFF 0x80040008L
#define OLE_E_CANT_GETMONIKER 0x80040009L
#define OLE_E_CANT_BINDTOSOURCE 0x8004000AL
#define OLE_E_STATIC 0x8004000BL
#define OLE_E_PROMPTSAVECANCELLED 0x8004000CL
#define OLE_E_INVALIDRECT 0x8004000DL
#define OLE_E_WRONGCOMPOBJ 0x8004000EL
#define OLE_E_INVALIDHWND 0x8004000FL
#define OLE_E_NOT_INPLACEACTIVE 0x80040010L
#define OLE_E_CANTCONVERT 0x80040011L
#define OLE_E_NOSTORAGE 0x80040012L
#define DV_E_FORMATETC 0x80040064L
#define DV_E_DVTARGETDEVICE 0x80040065L
#define DV_E_STGMEDIUM 0x80040066L
#define DV_E_STATDATA 0x80040067L
#define DV_E_LINDEX 0x80040068L
#define DV_E_TYMED 0x80040069L
#define DV_E_CLIPFORMAT 0x8004006AL
#define DV_E_DVASPECT 0x8004006BL
#define DV_E_DVTARGETDEVICE_SIZE 0x8004006CL
#define DV_E_NOIVIEWOBJECT 0x8004006DL
#define DRAGDROP_E_FIRST 0x80040100L
#define DRAGDROP_E_LAST 0x8004010FL
#define DRAGDROP_S_FIRST 0x00040100L
#define DRAGDROP_S_LAST 0x0004010FL
#define DRAGDROP_E_NOTREGISTERED 0x80040100L
#define DRAGDROP_E_ALREADYREGISTERED 0x80040101L
#define DRAGDROP_E_INVALIDHWND 0x80040102L
#define CLASSFACTORY_E_FIRST 0x80040110L
#define CLASSFACTORY_E_LAST 0x8004011FL
#define CLASSFACTORY_S_FIRST 0x00040110L
#define CLASSFACTORY_S_LAST 0x0004011FL
#define CLASS_E_NOAGGREGATION 0x80040110L
#define CLASS_E_CLASSNOTAVAILABLE 0x80040111L
#define MARSHAL_E_FIRST 0x80040120L
#define MARSHAL_E_LAST 0x8004012FL
#define MARSHAL_S_FIRST 0x00040120L
#define MARSHAL_S_LAST 0x0004012FL
#define DATA_E_FIRST 0x80040130L
#define DATA_E_LAST 0x8004013FL
#define DATA_S_FIRST 0x00040130L
#define DATA_S_LAST 0x0004013FL
#define VIEW_E_FIRST 0x80040140L
#define VIEW_E_LAST 0x8004014FL
#define VIEW_S_FIRST 0x00040140L
#define VIEW_S_LAST 0x0004014FL
#define VIEW_E_DRAW 0x80040140L
#define REGDB_E_FIRST 0x80040150L
#define REGDB_E_LAST 0x8004015FL
#define REGDB_S_FIRST 0x00040150L
#define REGDB_S_LAST 0x0004015FL
#define REGDB_E_READREGDB 0x80040150L
#define REGDB_E_WRITEREGDB 0x80040151L
#define REGDB_E_KEYMISSING 0x80040152L
#define REGDB_E_INVALIDVALUE 0x80040153L
#define REGDB_E_CLASSNOTREG 0x80040154L
#define REGDB_E_IIDNOTREG 0x80040155L
#define CACHE_E_FIRST 0x80040170L
#define CACHE_E_LAST 0x8004017FL
#define CACHE_S_FIRST 0x00040170L
#define CACHE_S_LAST 0x0004017FL
#define CACHE_E_NOCACHE_UPDATED 0x80040170L
#define OLEOBJ_E_FIRST 0x80040180L
#define OLEOBJ_E_LAST 0x8004018FL
#define OLEOBJ_S_FIRST 0x00040180L
#define OLEOBJ_S_LAST 0x0004018FL
#define OLEOBJ_E_NOVERBS 0x80040180L
#define OLEOBJ_E_INVALIDVERB 0x80040181L
#define CLIENTSITE_E_FIRST 0x80040190L
#define CLIENTSITE_E_LAST 0x8004019FL
#define CLIENTSITE_S_FIRST 0x00040190L
#define CLIENTSITE_S_LAST 0x0004019FL
#define INPLACE_E_NOTUNDOABLE 0x800401A0L
#define INPLACE_E_NOTOOLSPACE 0x800401A1L
#define INPLACE_E_FIRST 0x800401A0L
#define INPLACE_E_LAST 0x800401AFL
#define INPLACE_S_FIRST 0x000401A0L
#define INPLACE_S_LAST 0x000401AFL
#define ENUM_E_FIRST 0x800401B0L
#define ENUM_E_LAST 0x800401BFL
#define ENUM_S_FIRST 0x000401B0L
#define ENUM_S_LAST 0x000401BFL
#define CONVERT10_E_FIRST 0x800401C0L
#define CONVERT10_E_LAST 0x800401CFL
#define CONVERT10_S_FIRST 0x000401C0L
#define CONVERT10_S_LAST 0x000401CFL
#define CONVERT10_E_OLESTREAM_GET 0x800401C0L
#define CONVERT10_E_OLESTREAM_PUT 0x800401C1L
#define CONVERT10_E_OLESTREAM_FMT 0x800401C2L
#define CONVERT10_E_OLESTREAM_BITMAP_TO_DIB 0x800401C3L
#define CONVERT10_E_STG_FMT 0x800401C4L
#define CONVERT10_E_STG_NO_STD_STREAM 0x800401C5L
#define CONVERT10_E_STG_DIB_TO_BITMAP 0x800401C6L
#define CLIPBRD_E_FIRST 0x800401D0L
#define CLIPBRD_E_LAST 0x800401DFL
#define CLIPBRD_S_FIRST 0x000401D0L
#define CLIPBRD_S_LAST 0x000401DFL
#define CLIPBRD_E_CANT_OPEN 0x800401D0L
#define CLIPBRD_E_CANT_EMPTY 0x800401D1L
#define CLIPBRD_E_CANT_SET 0x800401D2L
#define CLIPBRD_E_BAD_DATA 0x800401D3L
#define CLIPBRD_E_CANT_CLOSE 0x800401D4L
#define MK_E_FIRST 0x800401E0L
#define MK_E_LAST 0x800401EFL
#define MK_S_FIRST 0x000401E0L
#define MK_S_LAST 0x000401EFL
#define MK_E_CONNECTMANUALLY 0x800401E0L
#define MK_E_EXCEEDEDDEADLINE 0x800401E1L
#define MK_E_NEEDGENERIC 0x800401E2L
#define MK_E_UNAVAILABLE 0x800401E3L
#define MK_E_SYNTAX 0x800401E4L
#define MK_E_NOOBJECT 0x800401E5L
#define MK_E_INVALIDEXTENSION 0x800401E6L
#define MK_E_INTERMEDIATEINTERFACENOTSUPPORTED 0x800401E7L
#define MK_E_NOTBINDABLE 0x800401E8L
#define MK_E_NOTBOUND 0x800401E9L
#define MK_E_CANTOPENFILE 0x800401EAL
#define MK_E_MUSTBOTHERUSER 0x800401EBL
#define MK_E_NOINVERSE 0x800401ECL
#define MK_E_NOSTORAGE 0x800401EDL
#define MK_E_NOPREFIX 0x800401EEL
#define MK_E_ENUMERATION_FAILED 0x800401EFL
#define CO_E_FIRST 0x800401F0L
#define CO_E_LAST 0x800401FFL
#define CO_S_FIRST 0x000401F0L
#define CO_S_LAST 0x000401FFL
#define CO_E_NOTINITIALIZED 0x800401F0L
#define CO_E_ALREADYINITIALIZED 0x800401F1L
#define CO_E_CANTDETERMINECLASS 0x800401F2L
#define CO_E_CLASSSTRING 0x800401F3L
#define CO_E_IIDSTRING 0x800401F4L
#define CO_E_APPNOTFOUND 0x800401F5L
#define CO_E_APPSINGLEUSE 0x800401F6L
#define CO_E_ERRORINAPP 0x800401F7L
#define CO_E_DLLNOTFOUND 0x800401F8L
#define CO_E_ERRORINDLL 0x800401F9L
#define CO_E_WRONGOSFORAPP 0x800401FAL
#define CO_E_OBJNOTREG 0x800401FBL
#define CO_E_OBJISREG 0x800401FCL
#define CO_E_OBJNOTCONNECTED 0x800401FDL
#define CO_E_APPDIDNTREG 0x800401FEL
#define CO_E_RELEASED 0x800401FFL
#define OLE_S_USEREG 0x00040000L
#define OLE_S_STATIC 0x00040001L
#define OLE_S_MAC_CLIPFORMAT 0x00040002L
#define DRAGDROP_S_DROP 0x00040100L
#define DRAGDROP_S_CANCEL 0x00040101L
#define DRAGDROP_S_USEDEFAULTCURSORS 0x00040102L
#define DATA_S_SAMEFORMATETC 0x00040130L
#define VIEW_S_ALREADY_FROZEN 0x00040140L
#define CACHE_S_FORMATETC_NOTSUPPORTED 0x00040170L
#define CACHE_S_SAMECACHE 0x00040171L
#define CACHE_S_SOMECACHES_NOTUPDATED 0x00040172L
#define OLEOBJ_S_INVALIDVERB 0x00040180L
#define OLEOBJ_S_CANNOT_DOVERB_NOW 0x00040181L
#define OLEOBJ_S_INVALIDHWND 0x00040182L
#define INPLACE_S_TRUNCATED 0x000401A0L
#define CONVERT10_S_NO_PRESENTATION 0x000401C0L
#define MK_S_REDUCED_TO_SELF 0x000401E2L
#define MK_S_ME 0x000401E4L
#define MK_S_HIM 0x000401E5L
#define MK_S_US 0x000401E6L
#define MK_S_MONIKERALREADYREGISTERED 0x000401E7L
#define CO_E_CLASS_CREATE_FAILED 0x80080001L
#define CO_E_SCM_ERROR 0x80080002L
#define CO_E_SCM_RPC_FAILURE 0x80080003L
#define CO_E_BAD_PATH 0x80080004L
#define CO_E_SERVER_EXEC_FAILURE 0x80080005L
#define CO_E_OBJSRV_RPC_FAILURE 0x80080006L
#define MK_E_NO_NORMALIZED 0x80080007L
#define CO_E_SERVER_STOPPING 0x80080008L
#define MEM_E_INVALID_ROOT 0x80080009L
#define MEM_E_INVALID_LINK 0x80080010L
#define MEM_E_INVALID_SIZE 0x80080011L
#define DISP_E_UNKNOWNINTERFACE 0x80020001L
#define DISP_E_MEMBERNOTFOUND 0x80020003L
#define DISP_E_PARAMNOTFOUND 0x80020004L
#define DISP_E_TYPEMISMATCH 0x80020005L
#define DISP_E_UNKNOWNNAME 0x80020006L
#define DISP_E_NONAMEDARGS 0x80020007L
#define DISP_E_BADVARTYPE 0x80020008L
#define DISP_E_EXCEPTION 0x80020009L
#define DISP_E_OVERFLOW 0x8002000AL
#define DISP_E_BADINDEX 0x8002000BL
#define DISP_E_UNKNOWNLCID 0x8002000CL
#define DISP_E_ARRAYISLOCKED 0x8002000DL
#define DISP_E_BADPARAMCOUNT 0x8002000EL
#define DISP_E_PARAMNOTOPTIONAL 0x8002000FL
#define DISP_E_BADCALLEE 0x80020010L
#define DISP_E_NOTACOLLECTION 0x80020011L
#define TYPE_E_BUFFERTOOSMALL 0x80028016L
#define TYPE_E_INVDATAREAD 0x80028018L
#define TYPE_E_UNSUPFORMAT 0x80028019L
#define TYPE_E_REGISTRYACCESS 0x8002801CL
#define TYPE_E_LIBNOTREGISTERED 0x8002801DL
#define TYPE_E_UNDEFINEDTYPE 0x80028027L
#define TYPE_E_QUALIFIEDNAMEDISALLOWED 0x80028028L
#define TYPE_E_INVALIDSTATE 0x80028029L
#define TYPE_E_WRONGTYPEKIND 0x8002802AL
#define TYPE_E_ELEMENTNOTFOUND 0x8002802BL
#define TYPE_E_AMBIGUOUSNAME 0x8002802CL
#define TYPE_E_NAMECONFLICT 0x8002802DL
#define TYPE_E_UNKNOWNLCID 0x8002802EL
#define TYPE_E_DLLFUNCTIONNOTFOUND 0x8002802FL
#define TYPE_E_BADMODULEKIND 0x800288BDL
#define TYPE_E_SIZETOOBIG 0x800288C5L
#define TYPE_E_DUPLICATEID 0x800288C6L
#define TYPE_E_INVALIDID 0x800288CFL
#define TYPE_E_TYPEMISMATCH 0x80028CA0L
#define TYPE_E_OUTOFBOUNDS 0x80028CA1L
#define TYPE_E_IOERROR 0x80028CA2L
#define TYPE_E_CANTCREATETMPFILE 0x80028CA3L
#define TYPE_E_CANTLOADLIBRARY 0x80029C4AL
#define TYPE_E_INCONSISTENTPROPFUNCS 0x80029C83L
#define TYPE_E_CIRCULARTYPE 0x80029C84L
#define STG_E_INVALIDFUNCTION 0x80030001L
#define STG_E_FILENOTFOUND 0x80030002L
#define STG_E_PATHNOTFOUND 0x80030003L
#define STG_E_TOOMANYOPENFILES 0x80030004L
#define STG_E_ACCESSDENIED 0x80030005L
#define STG_E_INVALIDHANDLE 0x80030006L
#define STG_E_INSUFFICIENTMEMORY 0x80030008L
#define STG_E_INVALIDPOINTER 0x80030009L
#define STG_E_NOMOREFILES 0x80030012L
#define STG_E_DISKISWRITEPROTECTED 0x80030013L
#define STG_E_SEEKERROR 0x80030019L
#define STG_E_WRITEFAULT 0x8003001DL
#define STG_E_READFAULT 0x8003001EL
#define STG_E_SHAREVIOLATION 0x80030020L
#define STG_E_LOCKVIOLATION 0x80030021L
#define STG_E_FILEALREADYEXISTS 0x80030050L
#define STG_E_INVALIDPARAMETER 0x80030057L
#define STG_E_MEDIUMFULL 0x80030070L
#define STG_E_ABNORMALAPIEXIT 0x800300FAL
#define STG_E_INVALIDHEADER 0x800300FBL
#define STG_E_INVALIDNAME 0x800300FCL
#define STG_E_UNKNOWN 0x800300FDL
#define STG_E_UNIMPLEMENTEDFUNCTION 0x800300FEL
#define STG_E_INVALIDFLAG 0x800300FFL
#define STG_E_INUSE 0x80030100L
#define STG_E_NOTCURRENT 0x80030101L
#define STG_E_REVERTED 0x80030102L
#define STG_E_CANTSAVE 0x80030103L
#define STG_E_OLDFORMAT 0x80030104L
#define STG_E_OLDDLL 0x80030105L
#define STG_E_SHAREREQUIRED 0x80030106L
#define STG_E_NOTFILEBASEDSTORAGE 0x80030107L
#define STG_E_EXTANTMARSHALLINGS 0x80030108L
#define STG_S_CONVERTED 0x00030200L
#define RPC_E_CALL_REJECTED 0x80010001L
#define RPC_E_CALL_CANCELED 0x80010002L
#define RPC_E_CANTPOST_INSENDCALL 0x80010003L
#define RPC_E_CANTCALLOUT_INASYNCCALL 0x80010004L
#define RPC_E_CANTCALLOUT_INEXTERNALCALL 0x80010005L
#define RPC_E_CONNECTION_TERMINATED 0x80010006L
#define RPC_E_SERVER_DIED 0x80010007L
#define RPC_E_CLIENT_DIED 0x80010008L
#define RPC_E_INVALID_DATAPACKET 0x80010009L
#define RPC_E_CANTTRANSMIT_CALL 0x8001000AL
#define RPC_E_CLIENT_CANTMARSHAL_DATA 0x8001000BL
#define RPC_E_CLIENT_CANTUNMARSHAL_DATA 0x8001000CL
#define RPC_E_SERVER_CANTMARSHAL_DATA 0x8001000DL
#define RPC_E_SERVER_CANTUNMARSHAL_DATA 0x8001000EL
#define RPC_E_INVALID_DATA 0x8001000FL
#define RPC_E_INVALID_PARAMETER 0x80010010L
#define RPC_E_CANTCALLOUT_AGAIN 0x80010011L
#define RPC_E_SERVER_DIED_DNE 0x80010012L
#define RPC_E_SYS_CALL_FAILED 0x80010100L
#define RPC_E_OUT_OF_RESOURCES 0x80010101L
#define RPC_E_ATTEMPTED_MULTITHREAD 0x80010102L
#define RPC_E_NOT_REGISTERED 0x80010103L
#define RPC_E_FAULT 0x80010104L
#define RPC_E_SERVERFAULT 0x80010105L
#define RPC_E_CHANGED_MODE 0x80010106L
#define RPC_E_INVALIDMETHOD 0x80010107L
#define RPC_E_DISCONNECTED 0x80010108L
#define RPC_E_RETRY 0x80010109L
#define RPC_E_SERVERCALL_RETRYLATER 0x8001010AL
#define RPC_E_SERVERCALL_REJECTED 0x8001010BL
#define RPC_E_INVALID_CALLDATA 0x8001010CL
#define RPC_E_CANTCALLOUT_ININPUTSYNCCALL 0x8001010DL
#define RPC_E_WRONG_THREAD 0x8001010EL
#define RPC_E_THREAD_NOT_INIT 0x8001010FL
#define RPC_E_UNEXPECTED 0x8001FFFFL
#define R2_BLACK 1
#define R2_NOTMERGEPEN 2
#define R2_MASKNOTPEN 3
#define R2_NOTCOPYPEN 4
#define R2_MASKPENNOT 5
#define R2_NOT 6
#define R2_XORPEN 7
#define R2_NOTMASKPEN 8
#define R2_MASKPEN 9
#define R2_NOTXORPEN 10
#define R2_NOP 11
#define R2_MERGENOTPEN 12 
#define R2_COPYPEN 13 
#define R2_MERGEPENNOT 14 
#define R2_MERGEPEN 15 
#define R2_WHITE 16 
#define R2_LAST 16
#define SRCCOPY 0x00CC0020U 
#define SRCPAINT 0x00EE0086U 
#define SRCAND 0x008800C6U 
#define SRCINVERT 0x00660046U 
#define SRCERASE 0x00440328U 
#define NOTSRCCOPY 0x00330008U 
#define NOTSRCERASE 0x001100A6U 
#define MERGECOPY 0x00C000CAU 
#define MERGEPAINT 0x00BB0226U 
#define PATCOPY 0x00F00021U 
#define PATPAINT 0x00FB0A09U 
#define PATINVERT 0x005A0049U 
#define DSTINVERT 0x00550009U 
#define BLACKNESS 0x00000042U 
#define WHITENESS 0x00FF0062U 
#define NOMIRRORBITMAP 0x80000000U 
#define CAPTUREBLT 0x40000000U 
#define GDI_ERROR 0xFFFFFFFFL
#define HGDI_ERROR DWORD(_cast,0xFFFFFFFFL)
#define NULLREGION 1
#define SIMPLEREGION 2
#define COMPLEXREGION 3
#define RGN_ERROR 0
#define RGN_AND 1
#define RGN_OR 2
#define RGN_XOR 3
#define RGN_DIFF 4
#define RGN_COPY 5
#define RGN_MIN RGN_AND
#define RGN_MAX RGN_COPY
#define BLACKONWHITE 1
#define WHITEONBLACK 2
#define COLORONCOLOR 3
#define HALFTONE 4
#define MAXSTRETCHBLTMODE 4
#define STRETCH_ANDSCANS BLACKONWHITE
#define STRETCH_ORSCANS WHITEONBLACK
#define STRETCH_DELETESCANS COLORONCOLOR
#define STRETCH_HALFTONE HALFTONE
#define ALTERNATE 1
#define WINDING 2
#define POLYFILL_LAST 2
#define LAYOUT_RTL 0x00000001
#define LAYOUT_BTT 0x00000002
#define LAYOUT_VBH 0x00000004
#define LAYOUT_ORIENTATIONMASK (LAYOUT_RTL | LAYOUT_BTT | LAYOUT_VBH)
#define LAYOUT_BITMAPORIENTATIONPRESERVED 0x00000008
#define TA_NOUPDATECP 0
#define TA_UPDATECP 1
#define TA_LEFT 0
#define TA_RIGHT 2
#define TA_CENTER 6
#define TA_TOP 0
#define TA_BOTTOM 8
#define TA_BASELINE 24
#define TA_RTLREADING 256
#define TA_MASK (TA_BASELINE+TA_CENTER+TA_UPDATECP+TA_RTLREADING)
#define VTA_BASELINE TA_BASELINE
#define VTA_LEFT TA_BOTTOM
#define VTA_RIGHT TA_TOP
#define VTA_CENTER TA_CENTER
#define VTA_BOTTOM TA_RIGHT
#define VTA_TOP TA_LEFT
#define ETO_OPAQUE 0x0002
#define ETO_CLIPPED 0x0004
#define ETO_GLYPH_INDEX 0x0010
#define ETO_RTLREADING 0x0080
#define ETO_NUMERICSLOCAL 0x0400
#define ETO_NUMERICSLATIN 0x0800
#define ETO_IGNORELANGUAGE 0x1000
#define ETO_PDY 0x2000
#define ASPECT_FILTERING 0x0001
#define DCB_RESET 0x0001
#define DCB_ACCUMULATE 0x0002
#define DCB_DIRTY DCB_ACCUMULATE
#define DCB_SET 0X0003
#define DCB_ENABLE 0x0004
#define DCB_DISABLE 0x0008
#define META_SETBKCOLOR 0x0201
#define META_SETBKMODE 0x0102
#define META_SETMAPMODE 0x0103
#define META_SETROP2 0x0104
#define META_SETRELABS 0x0105
#define META_SETPOLYFILLMODE 0x0106
#define META_SETSTRETCHBLTMODE 0x0107
#define META_SETTEXTCHAREXTRA 0x0108
#define META_SETTEXTCOLOR 0x0209
#define META_SETTEXTJUSTIFICATION 0x020A
#define META_SETWINDOWORG 0x020B
#define META_SETWINDOWEXT 0x020C
#define META_SETVIEWPORTORG 0x020D
#define META_SETVIEWPORTEXT 0x020E
#define META_OFFSETWINDOWORG 0x020F
#define META_SCALEWINDOWEXT 0x0410
#define META_OFFSETVIEWPORTORG 0x0211
#define META_SCALEVIEWPORTEXT 0x0412
#define META_LINETO 0x0213
#define META_MOVETO 0x0214
#define META_EXCLUDECLIPRECT 0x0415
#define META_INTERSECTCLIPRECT 0x0416
#define META_ARC 0x0817
#define META_ELLIPSE 0x0418
#define META_FLOODFILL 0x0419
#define META_PIE 0x081A
#define META_RECTANGLE 0x041B
#define META_ROUNDRECT 0x061C
#define META_PATBLT 0x061D
#define META_SAVEDC 0x001E
#define META_SETPIXEL 0x041F
#define META_OFFSETCLIPRGN 0x0220
#define META_TEXTOUT 0x0521
#define META_BITBLT 0x0922
#define META_STRETCHBLT 0x0B23
#define META_POLYGON 0x0324
#define META_POLYLINE 0x0325
#define META_ESCAPE 0x0626
#define META_RESTOREDC 0x0127
#define META_FILLREGION 0x0228
#define META_FRAMEREGION 0x0429
#define META_INVERTREGION 0x012A
#define META_PAINTREGION 0x012B
#define META_SELECTCLIPREGION 0x012C
#define META_SELECTOBJECT 0x012D
#define META_SETTEXTALIGN 0x012E
#define META_CHORD 0x0830
#define META_SETMAPPERFLAGS 0x0231
#define META_EXTTEXTOUT 0x0a32
#define META_SETDIBTODEV 0x0d33
#define META_SELECTPALETTE 0x0234
#define META_REALIZEPALETTE 0x0035
#define META_ANIMATEPALETTE 0x0436
#define META_SETPALENTRIES 0x0037
#define META_POLYPOLYGON 0x0538
#define META_RESIZEPALETTE 0x0139
#define META_DIBBITBLT 0x0940
#define META_DIBSTRETCHBLT 0x0b41
#define META_DIBCREATEPATTERNBRUSH 0x0142
#define META_STRETCHDIB 0x0f43
#define META_EXTFLOODFILL 0x0548
#define META_SETLAYOUT 0x0149
#define META_DELETEOBJECT 0x01f0
#define META_CREATEPALETTE 0x00f7
#define META_CREATEPATTERNBRUSH 0x01F9
#define META_CREATEPENINDIRECT 0x02FA
#define META_CREATEFONTINDIRECT 0x02FB
#define META_CREATEBRUSHINDIRECT 0x02FC
#define META_CREATEREGION 0x06FF
#define NEWFRAME 1
#define ABORTDOC_ 2
#define NEXTBAND 3
#define SETCOLORTABLE 4
#define GETCOLORTABLE 5
#define FLUSHOUTPUT 6
#define DRAFTMODE 7
#define QUERYESCSUPPORT 8
#define SETABORTPROC_ 9
#define STARTDOC_ 10
#define ENDDOC_ 11
#define GETPHYSPAGESIZE 12
#define GETPRINTINGOFFSET 13
#define GETSCALINGFACTOR 14
#define MFCOMMENT 15
#define GETPENWIDTH 16
#define SETCOPYCOUNT 17
#define SELECTPAPERSOURCE 18
#define DEVICEDATA 19
#define PASSTHROUGH 19
#define GETTECHNOLGY 20
#define GETTECHNOLOGY 20
#define SETLINECAP 21
#define SETLINEJOIN 22
#define bSETMITERLIMIT 23
#define BANDINFO 24
#define DRAWPATTERNRECT 25
#define GETVECTORPENSIZE 26
#define GETVECTORBRUSHSIZE 27
#define ENABLEDUPLEX 28
#define GETSETPAPERBINS 29
#define GETSETPRINTORIENT 30
#define ENUMPAPERBINS 31
#define SETDIBSCALING 32
#define EPSPRINTING 33
#define ENUMPAPERMETRICS 34
#define GETSETPAPERMETRICS 35
#define POSTSCRIPT_DATA 37
#define POSTSCRIPT_IGNORE 38
#define MOUSETRAILS 39
#define GETDEVICEUNITS 42
#define GETEXTENDEDTEXTMETRICS 256
#define GETEXTENTTABLE 257
#define GETPAIRKERNTABLE 258
#define GETTRACKKERNTABLE 259
#define bEXTTEXTOUT 512
#define GETFACENAME 513
#define DOWNLOADFACE 514
#define ENABLERELATIVEWIDTHS 768
#define ENABLEPAIRKERNING 769
#define SETKERNTRACK 770
#define SETALLJUSTVALUES 771
#define SETCHARSET 772
#define _STRETCHBLT 2048
#define METAFILE_DRIVER 2049
#define GETSETSCREENPARAMS 3072
#define QUERYDIBSUPPORT 3073
#define BEGIN_PATH 4096
#define CLIP_TO_PATH 4097
#define END_PATH 4098
#define EXT_DEVICE_CAPS 4099
#define RESTORE_CTM 4100
#define SAVE_CTM 4101
#define SET_ARC_DIRECTION 4102
#define SET_BACKGROUND_COLOR 4103
#define SET_POLY_MODE 4104
#define SET_SCREEN_ANGLE 4105
#define SET_SPREAD 4106
#define TRANSFORM_CTM 4107
#define SET_CLIP_BOX 4108
#define SET_BOUNDS 4109
#define SET_MIRROR_MODE 4110
#define OPENCHANNEL 4110
#define DOWNLOADHEADER 4111
#define CLOSECHANNEL 4112
#define POSTSCRIPT_PASSTHROUGH 4115
#define ENCAPSULATED_POSTSCRIPT 4116
#define POSTSCRIPT_IDENTIFY 4117 
#define POSTSCRIPT_INJECTION 4118 
#define CHECKJPEGFORMAT 4119
#define CHECKPNGFORMAT 4120
#define GET_PS_FEATURESETTING 4121 
#define SPCLPASSTHROUGH2 4568 
#define PSIDENT_GDICENTRIC 0
#define PSIDENT_PSCENTRIC 1
#define PSPROTOCOL_ASCII 0
#define PSPROTOCOL_BCP 1
#define PSPROTOCOL_TBCP 2
#define PSPROTOCOL_BINARY 3
#define QDI_SETDIBITS 1
#define QDI_GETDIBITS 2
#define QDI_DIBTOSCREEN 4
#define QDI_STRETCHDIB 8
#define SP_NOTREPORTED 0x4000
#define SP_ERROR (-1)
#define SP_APPABORT (-2)
#define SP_USERABORT (-3)
#define SP_OUTOFDISK (-4)
#define SP_OUTOFMEMORY (-5)
#define PR_JOBSTATUS 0x0000
#define OBJ_PEN 1
#define OBJ_BRUSH 2
#define OBJ_DC 3
#define OBJ_METADC 4
#define OBJ_PAL 5
#define OBJ_FONT 6
#define OBJ_BITMAP 7
#define OBJ_REGION 8
#define OBJ_METAFILE 9
#define OBJ_MEMDC 10
#define OBJ_EXTPEN 11
#define OBJ_ENHMETADC 12
#define OBJ_ENHMETAFILE 13
#define MWT_IDENTITY 1
#define MWT_LEFTMULTIPLY 2
#define MWT_RIGHTMULTIPLY 3
#define MWT_MIN MWT_IDENTITY
#define MWT_MAX MWT_RIGHTMULTIPLY
#define LCS_CALIBRATED_RGB 0x00000000L
#define LCS_DEVICE_RGB 0x00000001L
#define LCS_DEVICE_CMYK 0x00000002L
#define LCS_GM_BUSINESS 0x00000001L
#define LCS_GM_GRAPHICS 0x00000002L
#define LCS_GM_IMAGES 0x00000004L
#define CM_OUT_OF_GAMUT 255
#define CM_IN_GAMUT 0
#define BI_RGB 0L
#define BI_RLE8 1L
#define BI_RLE4 2L
#define BI_BITFIELDS 3L
#define BI_JPEG 4L
#define BI_PNG 5L
#define TCI_SRCCHARSET 1
#define TCI_SRCCODEPAGE 2
#define TCI_SRCFONTSIG 3
#define TMPF_FIXED_PITCH 0x01
#define TMPF_VECTOR 0x02
#define TMPF_DEVICE 0x08
#define TMPF_TRUETYPE 0x04
#define NTM_REGULAR 0x00000040L
#define NTM_BOLD 0x00000020L
#define NTM_ITALIC 0x00000001L
#define NTM_NONNEGATIVE_AC 0x00010000
#define NTM_PS_OPENTYPE 0x00020000
#define NTM_TT_OPENTYPE 0x00040000
#define NTM_MULTIPLEMASTER 0x00080000
#define NTM_TYPE1 0x00100000
#define NTM_DSIG 0x00200000
#define LF_FACESIZE 32
#define LF_FULLFACESIZE 64
#define OUT_DEFAULT_PRECIS 0
#define OUT_STRING_PRECIS 1
#define OUT_CHARACTER_PRECIS 2
#define OUT_STROKE_PRECIS 3
#define OUT_TT_PRECIS 4
#define OUT_DEVICE_PRECIS 5
#define OUT_RASTER_PRECIS 6
#define OUT_TT_ONLY_PRECIS 7
#define OUT_OUTLINE_PRECIS 8
#define OUT_SCREEN_OUTLINE_PRECIS 9
#define OUT_PS_ONLY_PRECIS 10
#define CLIP_DEFAULT_PRECIS 0
#define CLIP_CHARACTER_PRECIS 1
#define CLIP_STROKE_PRECIS 2
#define CLIP_MASK 0xf
#define CLIP_LH_ANGLES (1<<4)
#define CLIP_TT_ALWAYS (2<<4)
#define CLIP_DFA_DISABLE (4<<4)
#define CLIP_EMBEDDED (8<<4)
#define DEFAULT_QUALITY 0
#define DRAFT_QUALITY 1
#define PROOF_QUALITY 2
#define NONANTIALIASED_QUALITY 3
#define ANTIALIASED_QUALITY 4
#define CLEARTYPE_QUALITY 5
#define CLEARTYPE_NATURAL_QUALITY 6
#define DEFAULT_PITCH 0
#define FIXED_PITCH 1
#define VARIABLE_PITCH 2
#define MONO_FONT 8
#define ANSI_CHARSET 0
#define DEFAULT_CHARSET 1
#define SYMBOL_CHARSET 2
#define SHIFTJIS_CHARSET 128
#define HANGEUL_CHARSET 129
#define HANGUL_CHARSET 129
#define GB2312_CHARSET 134
#define CHINESEBIG5_CHARSET 136
#define OEM_CHARSET 255
#define JOHAB_CHARSET 130
#define HEBREW_CHARSET 177
#define ARABIC_CHARSET 178
#define GREEK_CHARSET 161
#define TURKISH_CHARSET 162
#define VIETNAMESE_CHARSET 163
#define THAI_CHARSET 222
#define EASTEUROPE_CHARSET 238
#define RUSSIAN_CHARSET 204
#define MAC_CHARSET 77
#define BALTIC_CHARSET 186
#define FS_LATIN1 0x00000001L
#define FS_LATIN2 0x00000002L
#define FS_CYRILLIC 0x00000004L
#define FS_GREEK 0x00000008L
#define FS_TURKISH 0x00000010L
#define FS_HEBREW 0x00000020L
#define FS_ARABIC 0x00000040L
#define FS_BALTIC 0x00000080L
#define FS_VIETNAMESE 0x00000100L
#define FS_THAI 0x00010000L
#define FS_JISJAPAN 0x00020000L
#define FS_CHINESESIMP 0x00040000L
#define FS_WANSUNG 0x00080000L
#define FS_CHINESETRAD 0x00100000L
#define FS_JOHAB 0x00200000L
#define FS_SYMBOL 0x80000000L
#define FF_DONTCARE (0<<4)
#define FF_ROMAN (1<<4)
#define FF_SWISS (2<<4)
#define FF_MODERN (3<<4)
#define FF_SCRIPT (4<<4)
#define FF_DECORATIVE (5<<4)
#define FW_DONTCARE 0
#define FW_THIN 100
#define FW_EXTRALIGHT 200
#define FW_LIGHT 300
#define FW_NORMAL 400
#define FW_MEDIUM 500
#define FW_SEMIBOLD 600
#define FW_BOLD 700
#define FW_EXTRABOLD 800
#define FW_HEAVY 900
#define FW_ULTRALIGHT FW_EXTRALIGHT
#define FW_REGULAR FW_NORMAL
#define FW_DEMIBOLD FW_SEMIBOLD
#define FW_ULTRABOLD FW_EXTRABOLD
#define FW_BLACK FW_HEAVY
#define PANOSE_COUNT 10
#define PAN_FAMILYTYPE_INDEX 0
#define PAN_SERIFSTYLE_INDEX 1
#define PAN_WEIGHT_INDEX 2
#define PAN_PROPORTION_INDEX 3
#define PAN_CONTRAST_INDEX 4
#define PAN_STROKEVARIATION_INDEX 5
#define PAN_ARMSTYLE_INDEX 6
#define PAN_LETTERFORM_INDEX 7
#define PAN_MIDLINE_INDEX 8
#define PAN_XHEIGHT_INDEX 9
#define PAN_CULTURE_LATIN 0
#define PAN_ANY 0
#define PAN_NO_FIT 1
#define PAN_FAMILY_TEXT_DISPLAY 2
#define PAN_FAMILY_SCRIPT 3
#define PAN_FAMILY_DECORATIVE 4
#define PAN_FAMILY_PICTORIAL 5
#define PAN_SERIF_COVE 2
#define PAN_SERIF_OBTUSE_COVE 3
#define PAN_SERIF_SQUARE_COVE 4
#define PAN_SERIF_OBTUSE_SQUARE_COVE 5
#define PAN_SERIF_SQUARE 6
#define PAN_SERIF_THIN 7
#define PAN_SERIF_BONE 8
#define PAN_SERIF_EXAGGERATED 9
#define PAN_SERIF_TRIANGLE 10
#define PAN_SERIF_NORMAL_SANS 11
#define PAN_SERIF_OBTUSE_SANS 12
#define PAN_SERIF_PERP_SANS 13
#define PAN_SERIF_FLARED 14
#define PAN_SERIF_ROUNDED 15
#define PAN_WEIGHT_VERY_LIGHT 2
#define PAN_WEIGHT_LIGHT 3
#define PAN_WEIGHT_THIN 4
#define PAN_WEIGHT_BOOK 5
#define PAN_WEIGHT_MEDIUM 6
#define PAN_WEIGHT_DEMI 7
#define PAN_WEIGHT_BOLD 8
#define PAN_WEIGHT_HEAVY 9
#define PAN_WEIGHT_BLACK 10
#define PAN_WEIGHT_NORD 11
#define PAN_PROP_OLD_STYLE 2
#define PAN_PROP_MODERN 3
#define PAN_PROP_EVEN_WIDTH 4
#define PAN_PROP_EXPANDED 5
#define PAN_PROP_CONDENSED 6
#define PAN_PROP_VERY_EXPANDED 7
#define PAN_PROP_VERY_CONDENSED 8
#define PAN_PROP_MONOSPACED 9
#define PAN_CONTRAST_NONE 2
#define PAN_CONTRAST_VERY_LOW 3
#define PAN_CONTRAST_LOW 4
#define PAN_CONTRAST_MEDIUM_LOW 5
#define PAN_CONTRAST_MEDIUM 6
#define PAN_CONTRAST_MEDIUM_HIGH 7
#define PAN_CONTRAST_HIGH 8
#define PAN_CONTRAST_VERY_HIGH 9
#define PAN_STROKE_GRADUAL_DIAG 2
#define PAN_STROKE_GRADUAL_TRAN 3
#define PAN_STROKE_GRADUAL_VERT 4
#define PAN_STROKE_GRADUAL_HORZ 5
#define PAN_STROKE_RAPID_VERT 6
#define PAN_STROKE_RAPID_HORZ 7
#define PAN_STROKE_INSTANT_VERT 8
#define PAN_STRAIGHT_ARMS_HORZ 2
#define PAN_STRAIGHT_ARMS_WEDGE 3
#define PAN_STRAIGHT_ARMS_VERT 4
#define PAN_STRAIGHT_ARMS_SINGLE_SERIF 5
#define PAN_STRAIGHT_ARMS_DOUBLE_SERIF 6
#define PAN_BENT_ARMS_HORZ 7
#define PAN_BENT_ARMS_WEDGE 8
#define PAN_BENT_ARMS_VERT 9
#define PAN_BENT_ARMS_SINGLE_SERIF 10
#define PAN_BENT_ARMS_DOUBLE_SERIF 11
#define PAN_LETT_NORMAL_CONTACT 2
#define PAN_LETT_NORMAL_WEIGHTED 3
#define PAN_LETT_NORMAL_BOXED 4
#define PAN_LETT_NORMAL_FLATTENED 5
#define PAN_LETT_NORMAL_ROUNDED 6
#define PAN_LETT_NORMAL_OFF_CENTER 7
#define PAN_LETT_NORMAL_SQUARE 8
#define PAN_LETT_OBLIQUE_CONTACT 9
#define PAN_LETT_OBLIQUE_WEIGHTED 10
#define PAN_LETT_OBLIQUE_BOXED 11
#define PAN_LETT_OBLIQUE_FLATTENED 12
#define PAN_LETT_OBLIQUE_ROUNDED 13
#define PAN_LETT_OBLIQUE_OFF_CENTER 14
#define PAN_LETT_OBLIQUE_SQUARE 15
#define PAN_MIDLINE_STANDARD_TRIMMED 2
#define PAN_MIDLINE_STANDARD_POINTED 3
#define PAN_MIDLINE_STANDARD_SERIFED 4
#define PAN_MIDLINE_HIGH_TRIMMED 5
#define PAN_MIDLINE_HIGH_POINTED 6
#define PAN_MIDLINE_HIGH_SERIFED 7
#define PAN_MIDLINE_CONSTANT_TRIMMED 8
#define PAN_MIDLINE_CONSTANT_POINTED 9
#define PAN_MIDLINE_CONSTANT_SERIFED 10
#define PAN_MIDLINE_LOW_TRIMMED 11
#define PAN_MIDLINE_LOW_POINTED 12
#define PAN_MIDLINE_LOW_SERIFED 13
#define PAN_XHEIGHT_CONSTANT_SMALL 2
#define PAN_XHEIGHT_CONSTANT_STD 3
#define PAN_XHEIGHT_CONSTANT_LARGE 4
#define PAN_XHEIGHT_DUCKING_SMALL 5
#define PAN_XHEIGHT_DUCKING_STD 6
#define PAN_XHEIGHT_DUCKING_LARGE 7
#define ELF_VENDOR_SIZE 4
#define ELF_VERSION 0
#define ELF_CULTURE_LATIN 0
#define RASTER_FONTTYPE 0x0001
#define DEVICE_FONTTYPE 0x002
#define TRUETYPE_FONTTYPE 0x004
#define PC_RESERVED 0x01
#define PC_EXPLICIT 0x02
#define PC_NOCOLLAPSE 0x04
#define TRANSPARENT 1
#define OPAQUE 2
#define BKMODE_LAST 2
#define GM_COMPATIBLE 1
#define GM_ADVANCED 2
#define GM_LAST 2
#define PT_CLOSEFIGURE 0x01
#define PT_LINETO 0x02
#define PT_BEZIERTO 0x04
#define PT_MOVETO 0x06
#define MM_TEXT 1
#define MM_LOMETRIC 2
#define MM_HIMETRIC 3
#define MM_LOENGLISH 4
#define MM_HIENGLISH 5
#define MM_TWIPS 6
#define MM_ISOTROPIC 7
#define MM_ANISOTROPIC 8
#define MM_MIN MM_TEXT
#define MM_MAX MM_ANISOTROPIC
#define MM_MAX_FIXEDSCALE MM_TWIPS
#define ABSOLUTE 1
#define RELATIVE 2
#define WHITE_BRUSH 0
#define LTGRAY_BRUSH 1
#define GRAY_BRUSH 2
#define DKGRAY_BRUSH 3
#define BLACK_BRUSH 4
#define NULL_BRUSH 5
#define HOLLOW_BRUSH NULL_BRUSH
#define WHITE_PEN 6
#define BLACK_PEN 7
#define NULL_PEN 8
#define OEM_FIXED_FONT 10
#define ANSI_FIXED_FONT 11
#define ANSI_VAR_FONT 12
#define SYSTEM_FONT 13
#define DEVICE_DEFAULT_FONT 14
#define DEFAULT_PALETTE 15
#define SYSTEM_FIXED_FONT 16
#define DEFAULT_GUI_FONT 17
#define DC_BRUSH 18
#define DC_PEN 19
#define STOCK_LAST 19
#define CLR_INVALID 0xFFFFFFFF
#define BS_SOLID 0
#define BS_NULL 1
#define BS_HOLLOW BS_NULL
#define BS_HATCHED 2
#define BS_PATTERN 3
#define BS_INDEXED 4
#define BS_DIBPATTERN 5
#define BS_DIBPATTERNPT 6
#define BS_PATTERN8X8 7
#define BS_DIBPATTERN8X8 8
#define BS_MONOPATTERN 9
#define HS_HORIZONTAL 0
#define HS_VERTICAL 1
#define HS_FDIAGONAL 2
#define HS_BDIAGONAL 3
#define HS_CROSS 4
#define HS_DIAGCROSS 5
#define PS_SOLID 0
#define PS_DASH 1
#define PS_DOT 2
#define PS_DASHDOT 3
#define PS_DASHDOTDOT 4
#define PS_NULL 5
#define PS_INSIDEFRAME 6
#define PS_USERSTYLE 7
#define PS_ALTERNATE 8
#define PS_STYLE_MASK 0x0000000F
#define PS_ENDCAP_ROUND 0x00000000
#define PS_ENDCAP_SQUARE 0x00000100
#define PS_ENDCAP_FLAT 0x00000200
#define PS_ENDCAP_MASK 0x00000F00
#define PS_JOIN_ROUND 0x00000000
#define PS_JOIN_BEVEL 0x00001000
#define PS_JOIN_MITER 0x00002000
#define PS_JOIN_MASK 0x0000F000
#define PS_COSMETIC 0x00000000
#define PS_GEOMETRIC 0x00010000
#define PS_TYPE_MASK 0x000F0000
#define AD_COUNTERCLOCKWISE 1
#define AD_CLOCKWISE 2
#define DRIVERVERSION 0
#define TECHNOLOGY 2
#define HORZSIZE 4
#define VERTSIZE 6
#define HORZRES 8
#define VERTRES 10
#define BITSPIXEL 12
#define PLANES 14
#define NUMBRUSHES 16
#define NUMPENS 18
#define NUMMARKERS 20
#define NUMFONTS 22
#define NUMCOLORS 24
#define PDEVICESIZE 26
#define CURVECAPS 28
#define LINECAPS 30
#define POLYGONALCAPS 32
#define TEXTCAPS 34
#define CLIPCAPS 36
#define RASTERCAPS 38
#define ASPECTX 40
#define ASPECTY 42
#define ASPECTXY 44
#define LOGPIXELSX 88
#define LOGPIXELSY 90
#define SIZEPALETTE 104
#define NUMRESERVED 106
#define COLORRES 108
#define PHYSICALWIDTH 110
#define PHYSICALHEIGHT 111
#define PHYSICALOFFSETX 112
#define PHYSICALOFFSETY 113
#define SCALINGFACTORX 114
#define SCALINGFACTORY 115
#define VREFRESH 116
#define DESKTOPVERTRES 117
#define DESKTOPHORZRES 118
#define BLTALIGNMENT 119
#define SHADEBLENDCAPS 120 
#define COLORMGMTCAPS 121 
#define DT_PLOTTER 0
#define DT_RASDISPLAY 1
#define DT_RASPRINTER 2
#define DT_RASCAMERA 3
#define DT_CHARSTREAM 4
#define DT_METAFILE 5
#define DT_DISPFILE 6
#define CC_NONE 0
#define CC_CIRCLES 1
#define CC_PIE 2
#define CC_CHORD 4
#define CC_ELLIPSES 8
#define CC_WIDE 16
#define CC_STYLED 32
#define CC_WIDESTYLED 64
#define CC_INTERIORS 128
#define CC_ROUNDRECT 256
#define LC_NONE 0
#define LC_POLYLINE 2
#define LC_MARKER 4
#define LC_POLYMARKER 8
#define LC_WIDE 16
#define LC_STYLED 32
#define LC_WIDESTYLED 64
#define LC_INTERIORS 128
#define PC_NONE 0
#define PC_POLYGON 1
#define PC_RECTANGLE 2
#define PC_WINDPOLYGON 4
#define PC_TRAPEZOID 4
#define PC_SCANLINE 8
#define PC_WIDE 16
#define PC_STYLED 32
#define PC_WIDESTYLED 64
#define PC_INTERIORS 128
#define PC_POLYPOLYGON 256
#define PC_PATHS 512
#define CP_NONE 0
#define CP_RECTANGLE 1
#define CP_REGION 2
#define TC_OP_CHARACTER 0x00000001
#define TC_OP_STROKE 0x00000002
#define TC_CP_STROKE 0x00000004
#define TC_CR_90 0x00000008
#define TC_CR_ANY 0x00000010
#define TC_SF_X_YINDEP 0x00000020
#define TC_SA_DOUBLE 0x00000040
#define TC_SA_INTEGER 0x00000080
#define TC_SA_CONTIN 0x00000100
#define TC_EA_DOUBLE 0x00000200
#define TC_IA_ABLE 0x00000400
#define TC_UA_ABLE 0x00000800
#define TC_SO_ABLE 0x00001000
#define TC_RA_ABLE 0x00002000
#define TC_VA_ABLE 0x00004000
#define TC_RESERVED 0x00008000
#define TC_SCROLLBLT 0x00010000
#define RC_BITBLT 1
#define RC_BANDING 2
#define RC_SCALING 4
#define RC_BITMAP64 8
#define RC_GDI20_OUTPUT 0x0010
#define RC_GDI20_STATE 0x0020
#define RC_SAVEBITMAP 0x0040
#define RC_DI_BITMAP 0x0080
#define RC_PALETTE 0x0100
#define RC_DIBTODEV 0x0200
#define RC_BIGFONT 0x0400
#define RC_STRETCHBLT 0x0800
#define RC_FLOODFILL 0x1000
#define RC_STRETCHDIB 0x2000
#define RC_OP_DX_OUTPUT 0x4000
#define RC_DEVBITS 0x8000
#define SB_NONE 0x00000000
#define SB_CONST_ALPHA 0x00000001
#define SB_PIXEL_ALPHA 0x00000002
#define SB_PREMULT_ALPHA 0x00000004
#define SB_GRAD_RECT 0x00000010
#define SB_GRAD_TRI 0x00000020
#define CM_NONE 0x00000000
#define CM_DEVICE_ICM 0x00000001
#define CM_GAMMA_RAMP 0x00000002
#define CM_CMYK_COLOR 0x00000004
#define DIB_RGB_COLORS 0
#define DIB_PAL_COLORS 1
#define SYSPAL_ERROR 0
#define SYSPAL_STATIC 1
#define SYSPAL_NOSTATIC 2
#define SYSPAL_NOSTATIC256 3
#define CBM_INIT 0x04L
#define FLOODFILLBORDER 0
#define FLOODFILLSURFACE 1
#define CCHDEVICENAME 32
#define CCHFORMNAME 32
#define DM_SPECVERSION 0x0400
#define DM_ORIENTATION 0x00000001L
#define DM_PAPERSIZE 0x00000002L
#define DM_PAPERLENGTH 0x00000004L
#define DM_PAPERWIDTH 0x00000008L
#define DM_SCALE 0x00000010L
#define DM_POSITION 0x00000020L
#define DM_NUP 0x00000040L
#define DM_DISPLAYORIENTATION 0x00000080L
#define DM_DEFAULTSOURCE 0x00000200L
#define DM_PRINTQUALITY 0x00000400L
#define DM_COLOR 0x00000800L
#define DM_DUPLEX 0x00001000L
#define DM_YRESOLUTION 0x00002000L
#define DM_TTOPTION 0x00004000L
#define DM_FORMNAME 0x00010000L
#define DM_LOGPIXELS 0x00020000L
#define DM_BITSPERPEL 0x00040000L
#define DM_PELSWIDTH 0x00080000L
#define DM_PELSHEIGHT 0x00100000L
#define DM_DISPLAYFLAGS 0x00200000L
#define DM_DISPLAYFREQUENCY 0x00400000L
#define DM_ICMMETHOD 0x00800000L
#define DM_ICMINTENT 0x01000000L
#define DM_MEDIATYPE 0x02000000L
#define DM_DITHERTYPE 0x04000000L
#define DM_PANNINGWIDTH 0x08000000L
#define DM_PANNINGHEIGHT 0x10000000L
#define DM_DISPLAYFIXEDOUTPUT 0x20000000L
#define DMORIENT_PORTRAIT 1
#define DMORIENT_LANDSCAPE 2
#define DMPAPER_LETTER 1
#define DMPAPER_FIRST DMPAPER_LETTER
#define DMPAPER_LETTERSMALL 2
#define DMPAPER_TABLOID 3
#define DMPAPER_LEDGER 4
#define DMPAPER_LEGAL 5
#define DMPAPER_STATEMENT 6
#define DMPAPER_EXECUTIVE 7
#define DMPAPER_A3 8
#define DMPAPER_A4 9
#define DMPAPER_A4SMALL 10
#define DMPAPER_A5 11
#define DMPAPER_B4 12
#define DMPAPER_B5 13
#define DMPAPER_FOLIO 14
#define DMPAPER_QUARTO 15
#define DMPAPER_10X14 16
#define DMPAPER_11X17 17
#define DMPAPER_NOTE 18
#define DMPAPER_ENV_9 19
#define DMPAPER_ENV_10 20
#define DMPAPER_ENV_11 21
#define DMPAPER_ENV_12 22
#define DMPAPER_ENV_14 23
#define DMPAPER_CSHEET 24
#define DMPAPER_DSHEET 25
#define DMPAPER_ESHEET 26
#define DMPAPER_ENV_DL 27
#define DMPAPER_ENV_C5 28
#define DMPAPER_ENV_C3 29
#define DMPAPER_ENV_C4 30
#define DMPAPER_ENV_C6 31
#define DMPAPER_ENV_C65 32
#define DMPAPER_ENV_B4 33
#define DMPAPER_ENV_B5 34
#define DMPAPER_ENV_B6 35
#define DMPAPER_ENV_ITALY 36
#define DMPAPER_ENV_MONARCH 37
#define DMPAPER_ENV_PERSONAL 38
#define DMPAPER_FANFOLD_US 39
#define DMPAPER_FANFOLD_STD_GERMAN 40
#define DMPAPER_FANFOLD_LGL_GERMAN 41
#define DMPAPER_ISO_B4 42
#define DMPAPER_JAPANESE_POSTCARD 43
#define DMPAPER_9X11 44
#define DMPAPER_10X11 45
#define DMPAPER_15X11 46
#define DMPAPER_ENV_INVITE 47
#define DMPAPER_RESERVED_48 48
#define DMPAPER_RESERVED_49 49
#define DMPAPER_LETTER_EXTRA 50
#define DMPAPER_LEGAL_EXTRA 51
#define DMPAPER_TABLOID_EXTRA 52
#define DMPAPER_A4_EXTRA 53
#define DMPAPER_LETTER_TRANSVERSE 54
#define DMPAPER_A4_TRANSVERSE 55
#define DMPAPER_LETTER_EXTRA_TRANSVERSE 56
#define DMPAPER_A_PLUS 57
#define DMPAPER_B_PLUS 58
#define DMPAPER_LETTER_PLUS 59
#define DMPAPER_A4_PLUS 60
#define DMPAPER_A5_TRANSVERSE 61
#define DMPAPER_B5_TRANSVERSE 62
#define DMPAPER_A3_EXTRA 63
#define DMPAPER_A5_EXTRA 64
#define DMPAPER_B5_EXTRA 65
#define DMPAPER_A2 66
#define DMPAPER_A3_TRANSVERSE 67
#define DMPAPER_A3_EXTRA_TRANSVERSE 68
#define DMPAPER_DBL_JAPANESE_POSTCARD 69 
#define DMPAPER_A6 70 
#define DMPAPER_JENV_KAKU2 71 
#define DMPAPER_JENV_KAKU3 72 
#define DMPAPER_JENV_CHOU3 73 
#define DMPAPER_JENV_CHOU4 74 
#define DMPAPER_LETTER_ROTATED 75 
#define DMPAPER_A3_ROTATED 76 
#define DMPAPER_A4_ROTATED 77 
#define DMPAPER_A5_ROTATED 78 
#define DMPAPER_B4_JIS_ROTATED 79 
#define DMPAPER_B5_JIS_ROTATED 80 
#define DMPAPER_JAPANESE_POSTCARD_ROTATED 81 
#define DMPAPER_DBL_JAPANESE_POSTCARD_ROTATED 82 
#define DMPAPER_A6_ROTATED 83 
#define DMPAPER_JENV_KAKU2_ROTATED 84 
#define DMPAPER_JENV_KAKU3_ROTATED 85 
#define DMPAPER_JENV_CHOU3_ROTATED 86 
#define DMPAPER_JENV_CHOU4_ROTATED 87 
#define DMPAPER_B6_JIS 88 
#define DMPAPER_B6_JIS_ROTATED 89 
#define DMPAPER_12X11 90 
#define DMPAPER_JENV_YOU4 91 
#define DMPAPER_JENV_YOU4_ROTATED 92 
#define DMPAPER_P16K 93 
#define DMPAPER_P32K 94 
#define DMPAPER_P32KBIG 95 
#define DMPAPER_PENV_1 96 
#define DMPAPER_PENV_2 97 
#define DMPAPER_PENV_3 98 
#define DMPAPER_PENV_4 99 
#define DMPAPER_PENV_5 100 
#define DMPAPER_PENV_6 101 
#define DMPAPER_PENV_7 102 
#define DMPAPER_PENV_8 103 
#define DMPAPER_PENV_9 104 
#define DMPAPER_PENV_10 105 
#define DMPAPER_P16K_ROTATED 106 
#define DMPAPER_P32K_ROTATED 107 
#define DMPAPER_P32KBIG_ROTATED 108 
#define DMPAPER_PENV_1_ROTATED 109 
#define DMPAPER_PENV_2_ROTATED 110 
#define DMPAPER_PENV_3_ROTATED 111 
#define DMPAPER_PENV_4_ROTATED 112 
#define DMPAPER_PENV_5_ROTATED 113 
#define DMPAPER_PENV_6_ROTATED 114 
#define DMPAPER_PENV_7_ROTATED 115 
#define DMPAPER_PENV_8_ROTATED 116 
#define DMPAPER_PENV_9_ROTATED 117 
#define DMPAPER_PENV_10_ROTATED 118 
#define DMPAPER_LAST DMPAPER_PENV_10_ROTATED
#define DMPAPER_USER 256
#define DMBIN_UPPER 1
#define DMBIN_FIRST DMBIN_UPPER
#define DMBIN_ONLYONE 1
#define DMBIN_LOWER 2
#define DMBIN_MIDDLE 3
#define DMBIN_MANUAL 4
#define DMBIN_ENVELOPE 5
#define DMBIN_ENVMANUAL 6
#define DMBIN_AUTO 7
#define DMBIN_TRACTOR 8
#define DMBIN_SMALLFMT 9
#define DMBIN_LARGEFMT 10
#define DMBIN_LARGECAPACITY 11
#define DMBIN_CASSETTE 14
#define DMBIN_FORMSOURCE 15
#define DMBIN_LAST DMBIN_FORMSOURCE
#define DMBIN_USER 256
#define DMRES_DRAFT (-1)
#define DMRES_LOW (-2)
#define DMRES_MEDIUM (-3)
#define DMRES_HIGH (-4)
#define DMCOLOR_MONOCHROME 1
#define DMCOLOR_COLOR 2
#define DMDUP_SIMPLEX 1
#define DMDUP_VERTICAL 2
#define DMDUP_HORIZONTAL 3
#define DMTT_BITMAP 1
#define DMTT_DOWNLOAD 2
#define DMTT_SUBDEV 3
#define DMTT_DOWNLOAD_OUTLINE 4
#define DMCOLLATE_FALSE 0
#define DMCOLLATE_TRUE 1
#define DMDO_DEFAULT 0
#define DMDO_90 1
#define DMDO_180 2
#define DMDO_270 3
#define DMDFO_DEFAULT 0
#define DMDFO_STRETCH 1
#define DMDFO_CENTER 2
#define DM_GRAYSCALE 0x00000001
#define DM_INTERLACED 0x00000002
#define DMICMMETHOD_NONE 1
#define DMICMMETHOD_SYSTEM 2
#define DMICMMETHOD_DRIVER 3
#define DMICMMETHOD_DEVICE 4
#define DMICMMETHOD_USER 256
#define DMICM_SATURATE 1
#define DMICM_CONTRAST 2
#define DMICM_COLORMETRIC 3
#define DMICM_ABS_COLORIMETRIC 4 
#define DMICM_USER 256
#define DMMEDIA_STANDARD 1
#define DMMEDIA_TRANSPARENCY 2
#define DMMEDIA_GLOSSY 3
#define DMMEDIA_USER 256
#define DMDITHER_NONE 1
#define DMDITHER_COARSE 2
#define DMDITHER_FINE 3
#define DMDITHER_LINEART 4
#define DMDITHER_ERRORDIFFUSION 5
#define DMDITHER_RESERVED6 6
#define DMDITHER_RESERVED7 7
#define DMDITHER_RESERVED8 8
#define DMDITHER_RESERVED9 9
#define DMDITHER_GRAYSCALE 10
#define DMDITHER_USER 256
#define DISPLAY_DEVICE_ATTACHED_TO_DESKTOP 0x00000001
#define DISPLAY_DEVICE_MULTI_DRIVER 0x00000002
#define DISPLAY_DEVICE_PRIMARY_DEVICE 0x00000004
#define DISPLAY_DEVICE_MIRRORING_DRIVER 0x00000008
#define DISPLAY_DEVICE_VGA_COMPATIBLE 0x00000010
#define DISPLAY_DEVICE_REMOVABLE 0x00000020
#define DISPLAY_DEVICE_MODESPRUNED 0x08000000
#define DISPLAY_DEVICE_REMOTE 0x04000000
#define DISPLAY_DEVICE_DISCONNECT 0x02000000
#define DISPLAY_DEVICE_ACTIVE 0x00000001
#define DISPLAY_DEVICE_ATTACHED 0x00000002
#define RDH_RECTANGLES 1
#define GGO_METRICS 0
#define GGO_BITMAP 1
#define GGO_NATIVE 2
#define GGO_BEZIER 3
#define GGO_GRAY2_BITMAP 4
#define GGO_GRAY4_BITMAP 5
#define GGO_GRAY8_BITMAP 6
#define GGO_GLYPH_INDEX 0x0080
#define GGO_UNHINTED 0x0100
#define TT_POLYGON_TYPE 24
#define TT_PRIM_LINE 1
#define TT_PRIM_QSPLINE 2
#define TT_PRIM_CSPLINE 3
#define GCP_DBCS 0x0001
#define GCP_REORDER 0x0002
#define GCP_USEKERNING 0x0008
#define GCP_GLYPHSHAPE 0x0010
#define GCP_LIGATE 0x0020
#define GCP_DIACRITIC 0x0100
#define GCP_KASHIDA 0x0400
#define GCP_ERROR 0x8000
#define FLI_MASK 0x103B
#define GCP_JUSTIFY 0x00010000L
#define FLI_GLYPHS 0x00040000L
#define GCP_CLASSIN 0x00080000L
#define GCP_MAXEXTENT 0x00100000L
#define GCP_JUSTIFYIN 0x00200000L
#define GCP_DISPLAYZWG 0x00400000L
#define GCP_SYMSWAPOFF 0x00800000L
#define GCP_NUMERICOVERRIDE 0x01000000L
#define GCP_NEUTRALOVERRIDE 0x02000000L
#define GCP_NUMERICSLATIN 0x04000000L
#define GCP_NUMERICSLOCAL 0x08000000L
#define GCPCLASS_LATIN 1
#define GCPCLASS_HEBREW 2
#define GCPCLASS_ARABIC 2
#define GCPCLASS_NEUTRAL 3
#define GCPCLASS_LOCALNUMBER 4
#define GCPCLASS_LATINNUMBER 5
#define GCPCLASS_LATINNUMERICTERMINATOR 6
#define GCPCLASS_LATINNUMERICSEPARATOR 7
#define GCPCLASS_NUMERICSEPARATOR 8
#define GCPCLASS_PREBOUNDLTR 0x80
#define GCPCLASS_PREBOUNDRTL 0x40
#define GCPCLASS_POSTBOUNDLTR 0x20
#define GCPCLASS_POSTBOUNDRTL 0x10
#define GCPGLYPH_LINKBEFORE 0x8000
#define GCPGLYPH_LINKAFTER 0x4000
#define TT_AVAILABLE 0x0001
#define TT_ENABLED 0x0002
#define PFD_TYPE_RGBA 0
#define PFD_TYPE_COLORINDEX 1
#define PFD_MAIN_PLANE 0
#define PFD_OVERLAY_PLANE 1
#define PFD_UNDERLAY_PLANE (-1)
#define PFD_DOUBLEBUFFER 0x00000001
#define PFD_STEREO 0x00000002
#define PFD_DRAW_TO_WINDOW 0x00000004
#define PFD_DRAW_TO_BITMAP 0x00000008
#define PFD_SUPPORT_GDI 0x00000010
#define PFD_SUPPORT_OPENGL 0x00000020
#define PFD_GENERIC_FORMAT 0x00000040
#define PFD_NEED_PALETTE 0x00000080
#define PFD_NEED_SYSTEM_PALETTE 0x00000100
#define PFD_SWAP_EXCHANGE 0x00000200
#define PFD_SWAP_COPY 0x00000400
#define PFD_SWAP_LAYER_BUFFERS 0x00000800
#define PFD_GENERIC_ACCELERATED 0x00001000
#define PFD_SUPPORT_DIRECTDRAW 0x00002000
#define PFD_DEPTH_DONTCARE 0x20000000
#define PFD_DOUBLEBUFFER_DONTCARE 0x40000000
#define PFD_STEREO_DONTCARE 0x80000000
#define DM_UPDATE 1
#define DM_COPY 2
#define DM_PROMPT 4
#define DM_MODIFY 8
#define DM_IN_BUFFER DM_MODIFY
#define DM_IN_PROMPT DM_PROMPT
#define DM_OUT_BUFFER DM_COPY
#define DM_OUT_DEFAULT DM_UPDATE
#define DC_FIELDS 1
#define DC_PAPERS 2
#define DC_PAPERSIZE 3
#define DC_MINEXTENT 4
#define DC_MAXEXTENT 5
#define DC_BINS 6
#define DC_DUPLEX 7
#define DC_SIZE 8
#define DC_EXTRA 9
#define DC_VERSION 10
#define DC_DRIVER 11
#define DC_BINNAMES 12
#define DC_ENUMRESOLUTIONS 13
#define DC_FILEDEPENDENCIES 14
#define DC_TRUETYPE 15
#define DC_PAPERNAMES 16
#define DC_ORIENTATION 17
#define DC_COPIES 18
#define DC_BINADJUST 19
#define DC_EMF_COMPLIANT 20
#define DC_DATATYPE_PRODUCED 21
#define DC_COLLATE 22
#define DC_MANUFACTURER 23
#define DC_MODEL 24
#define DC_PERSONALITY 25
#define DC_PRINTRATE 26
#define DC_PRINTRATEUNIT 27
#define PRINTRATEUNIT_PPM 1
#define PRINTRATEUNIT_CPS 2
#define PRINTRATEUNIT_LPM 3
#define PRINTRATEUNIT_IPM 4
#define DC_PRINTERMEM 28
#define DC_MEDIAREADY 29
#define DC_STAPLE 30
#define DC_PRINTRATEPPM 31
#define DC_COLORDEVICE 32
#define DC_NUP 33
#define DC_MEDIATYPENAMES 34
#define DC_MEDIATYPES 35
#define DCTT_BITMAP 0x0000001L
#define DCTT_DOWNLOAD 0x0000002L
#define DCTT_SUBDEV 0x0000004L
#define DCTT_DOWNLOAD_OUTLINE 0x0000008L
#define DCBA_FACEUPNONE 0x0000
#define DCBA_FACEUPCENTER 0x0001
#define DCBA_FACEUPLEFT 0x0002
#define DCBA_FACEUPRIGHT 0x0003
#define DCBA_FACEDOWNNONE 0x0100
#define DCBA_FACEDOWNCENTER 0x0101
#define DCBA_FACEDOWNLEFT 0x0102
#define DCBA_FACEDOWNRIGHT 0x0103
#define CA_NEGATIVE 0x0001
#define CA_LOG_FILTER 0x0002
#define ILLUMINANT_DEVICE_DEFAULT 0
#define ILLUMINANT_A 1
#define ILLUMINANT_B 2
#define ILLUMINANT_C 3
#define ILLUMINANT_D50 4
#define ILLUMINANT_D55 5
#define ILLUMINANT_D65 6
#define ILLUMINANT_D75 7
#define ILLUMINANT_F2 8
#define ILLUMINANT_MAX_INDEX ILLUMINANT_F2
#define ILLUMINANT_TUNGSTEN ILLUMINANT_A
#define ILLUMINANT_DAYLIGHT ILLUMINANT_C
#define ILLUMINANT_FLUORESCENT ILLUMINANT_F2
#define ILLUMINANT_NTSC ILLUMINANT_C
#define RGB_GAMMA_MIN WORD(_cast,02500)
#define RGB_GAMMA_MAX WORD(_cast, 65000)
#define REFERENCE_WHITE_MIN WORD(_cast,6000)
#define REFERENCE_WHITE_MAX WORD(_cast,10000)
#define REFERENCE_BLACK_MIN WORD(_cast,0)
#define REFERENCE_BLACK_MAX WORD(_cast,4000)
#define COLOR_ADJ_MIN -100
#define DI_APPBANDING 0x0001
#define FONTMAPPER_MAX 10
#define ICM_OFF 1
#define ICM_ON 2
#define ICM_QUERY 3
#define ICM_DONE_OUTSIDEDC 4
#define ENHMETA_SIGNATURE 0x464D4520
#define ENHMETA_STOCK_OBJECT 0x80000000
#define EMR_HEADER 1
#define EMR_POLYBEZIER 2
#define EMR_POLYGON 3
#define EMR_POLYLINE 4
#define EMR_POLYBEZIERTO 5
#define EMR_POLYLINETO 6
#define EMR_POLYPOLYLINE 7
#define EMR_POLYPOLYGON 8
#define EMR_SETWINDOWEXTEX 9
#define EMR_SETWINDOWORGEX 10
#define EMR_SETVIEWPORTEXTEX 11
#define EMR_SETVIEWPORTORGEX 12
#define EMR_SETBRUSHORGEX 13
#define EMR_EOF 14
#define EMR_SETPIXELV 15
#define EMR_SETMAPPERFLAGS 16
#define EMR_SETMAPMODE 17
#define EMR_SETBKMODE 18
#define EMR_SETPOLYFILLMODE 19
#define EMR_SETROP2 20
#define EMR_SETSTRETCHBLTMODE 21
#define EMR_SETTEXTALIGN 22
#define EMR_SETCOLORADJUSTMENT 23
#define EMR_SETTEXTCOLOR 24
#define EMR_SETBKCOLOR 25
#define EMR_OFFSETCLIPRGN 26
#define EMR_MOVETOEX 27
#define EMR_SETMETARGN 28
#define EMR_EXCLUDECLIPRECT 29
#define EMR_INTERSECTCLIPRECT 30
#define EMR_SCALEVIEWPORTEXTEX 31
#define EMR_SCALEWINDOWEXTEX 32
#define EMR_SAVEDC 33
#define EMR_RESTOREDC 34
#define EMR_SETWORLDTRANSFORM 35
#define EMR_MODIFYWORLDTRANSFORM 36
#define EMR_SELECTOBJECT 37
#define EMR_CREATEPEN 38
#define EMR_CREATEBRUSHINDIRECT 39
#define EMR_DELETEOBJECT 40
#define EMR_ANGLEARC 41
#define EMR_ELLIPSE 42
#define EMR_RECTANGLE 43
#define EMR_ROUNDRECT 44
#define EMR_ARC 45
#define EMR_CHORD 46
#define EMR_PIE 47
#define EMR_SELECTPALETTE 48
#define EMR_CREATEPALETTE 49
#define EMR_SETPALETTEENTRIES 50
#define EMR_RESIZEPALETTE 51
#define EMR_REALIZEPALETTE 52
#define EMR_EXTFLOODFILL 53
#define EMR_LINETO 54
#define EMR_ARCTO 55
#define EMR_POLYDRAW 56
#define EMR_SETARCDIRECTION 57
#define EMR_SETMITERLIMIT 58
#define EMR_BEGINPATH 59
#define EMR_ENDPATH 60
#define EMR_CLOSEFIGURE 61
#define EMR_FILLPATH 62
#define EMR_STROKEANDFILLPATH 63
#define EMR_STROKEPATH 64
#define EMR_FLATTENPATH 65
#define EMR_WIDENPATH 66
#define EMR_SELECTCLIPPATH 67
#define EMR_ABORTPATH 68
#define EMR_GDICOMMENT 70
#define EMR_FILLRGN 71
#define EMR_FRAMERGN 72
#define EMR_INVERTRGN 73
#define EMR_PAINTRGN 74
#define EMR_EXTSELECTCLIPRGN 75
#define EMR_BITBLT 76
#define EMR_STRETCHBLT 77
#define EMR_MASKBLT 78
#define EMR_PLGBLT 79
#define EMR_SETDIBITSTODEVICE 80
#define EMR_STRETCHDIBITS 81
#define EMR_EXTCREATEFONTINDIRECTW 82
#define EMR_EXTTEXTOUTA 83
#define EMR_EXTTEXTOUTW 84
#define EMR_POLYBEZIER16 85
#define EMR_POLYGON16 86
#define EMR_POLYLINE16 87
#define EMR_POLYBEZIERTO16 88
#define EMR_POLYLINETO16 89
#define EMR_POLYPOLYLINE16 90
#define EMR_POLYPOLYGON16 91
#define EMR_POLYDRAW16 92
#define EMR_CREATEMONOBRUSH 93
#define EMR_CREATEDIBPATTERNBRUSHPT 94
#define EMR_EXTCREATEPEN 95
#define EMR_POLYTEXTOUTA 96
#define EMR_POLYTEXTOUTW 97
#define EMR_SETICMMODE 98
#define EMR_CREATECOLORSPACE 99
#define EMR_SETCOLORSPACE 100
#define EMR_DELETECOLORSPACE 101
#define EMR_GLSRECORD 102
#define EMR_GLSBOUNDEDRECORD 103
#define EMR_PIXELFORMAT 104
#define EMR_RESERVED_105 105
#define EMR_RESERVED_106 106
#define EMR_RESERVED_107 107
#define EMR_RESERVED_108 108
#define EMR_RESERVED_109 109
#define EMR_RESERVED_110 110
#define EMR_COLORCORRECTPALETTE 111
#define EMR_SETICMPROFILEA 112
#define EMR_SETICMPROFILEW 113
#define EMR_ALPHABLEND 114
#define EMR_SETLAYOUT 115
#define EMR_TRANSPARENTBLT 116
#define EMR_RESERVED_117 117
#define EMR_GRADIENTFILL 118
#define EMR_RESERVED_119 119
#define EMR_RESERVED_120 120
#define EMR_COLORMATCHTOTARGETW 121
#define EMR_CREATECOLORSPACEW 122
#define EMR_MIN 1
#define EMR_MAX 122
#define GDICOMMENT_IDENTIFIER 0x43494447
#define GDICOMMENT_WINDOWS_METAFILE 0x80000001
#define GDICOMMENT_BEGINGROUP 0x00000002
#define GDICOMMENT_ENDGROUP 0x00000003
#define GDICOMMENT_MULTIFORMATS 0x40000004
#define EPS_SIGNATURE 0x46535045
#define GDICOMMENT_UNICODE_STRING 0x00000040
#define GDICOMMENT_UNICODE_END 0x00000080
#define WGL_FONT_LINES 0
#define WGL_FONT_POLYGONS 1
#define COLOR_ADJ_MAX SHORTINT(_cast, 100)
#define INTERNET_INVALID_PORT_NUMBER 0
#define INTERNET_DEFAULT_FTP_PORT 21
#define INTERNET_DEFAULT_GOPHER_PORT 70
#define INTERNET_DEFAULT_HTTP_PORT 80
#define INTERNET_DEFAULT_HTTPS_PORT 443
#define INTERNET_DEFAULT_SOCKS_PORT 1080
#define MAX_CACHE_ENTRY_INFO_SIZE 4096
#define INTERNET_MAX_HOST_NAME_LENGTH 256
#define INTERNET_MAX_USER_NAME_LENGTH 128
#define INTERNET_MAX_PASSWORD_LENGTH 128
#define INTERNET_MAX_PORT_NUMBER_LENGTH 5
#define INTERNET_MAX_PORT_NUMBER_VALUE 65535
#define INTERNET_MAX_PATH_LENGTH 2048
#define INTERNET_MAX_PROTOCOL_NAME "gopher"
#define INTERNET_MAX_SCHEME_LENGTH 32
#define _INTERNET_MAX_URL_LENGTH INTERNET_MAX_SCHEME_LENGTH + 3 +INTERNET_MAX_PATH_LENGTH
#define INTERNET_KEEP_ALIVE_UNKNOWN 0xFFFFFFFF
#define INTERNET_KEEP_ALIVE_ENABLED 1
#define INTERNET_KEEP_ALIVE_DISABLED 0
#define INTERNET_REQFLAG_FROM_CACHE 0x00000001
#define INTERNET_REQFLAG_ASYNC 0x00000002
#define INTERNET_REQFLAG_VIA_PROXY 0x00000004
#define INTERNET_REQFLAG_NO_HEADERS 0x00000008
#define INTERNET_REQFLAG_PASSIVE 0x00000010
#define INTERNET_REQFLAG_CACHE_WRITE_DISABLED 0x00000040
#define INTERNET_REQFLAG_NET_TIMEOUT 0x00000080
#define INTERNET_FLAG_RELOAD 0x80000000
#define INTERNET_FLAG_RAW_DATA 0x40000000
#define INTERNET_FLAG_EXISTING_CONNECT 0x20000000
#define INTERNET_FLAG_ASYNC 0x10000000
#define INTERNET_FLAG_PASSIVE 0x08000000
#define INTERNET_FLAG_NO_CACHE_WRITE 0x04000000
#define INTERNET_FLAG_DONT_CACHE INTERNET_FLAG_NO_CACHE_WRITE
#define INTERNET_FLAG_MAKE_PERSISTENT 0x02000000
#define INTERNET_FLAG_FROM_CACHE 0x01000000
#define INTERNET_FLAG_OFFLINE INTERNET_FLAG_FROM_CACHE
#define INTERNET_FLAG_SECURE 0x00800000
#define INTERNET_FLAG_KEEP_CONNECTION 0x00400000
#define INTERNET_FLAG_NO_AUTO_REDIRECT 0x00200000
#define INTERNET_FLAG_READ_PREFETCH 0x00100000
#define INTERNET_FLAG_NO_COOKIES 0x00080000
#define INTERNET_FLAG_NO_AUTH 0x00040000
#define INTERNET_FLAG_RESTRICTED_ZONE 0x00020000
#define INTERNET_FLAG_CACHE_IF_NET_FAIL 0x00010000
#define INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTP 0x00008000
#define INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTPS 0x00004000
#define INTERNET_FLAG_IGNORE_CERT_DATE_INVALID 0x00002000
#define INTERNET_FLAG_IGNORE_CERT_CN_INVALID 0x00001000
#define INTERNET_FLAG_BGUPDATE 0x00000008
#define INTERNET_FLAG_MUST_CACHE_REQUEST 0x00000010
#define INTERNET_FLAG_RESYNCHRONIZE 0x00000800
#define INTERNET_FLAG_HYPERLINK 0x00000400
#define INTERNET_FLAG_NO_UI 0x00000200
#define INTERNET_FLAG_PRAGMA_NOCACHE 0x00000100
#define INTERNET_FLAG_CACHE_ASYNC 0x00000080
#define INTERNET_FLAG_FORMS_SUBMIT 0x00000040
#define INTERNET_FLAG_FWD_BACK 0x00000020
#define INTERNET_FLAG_NEED_FILE 0x00000010
#define FTP_TRANSFER_TYPE_ASCII 0x00000001
#define INTERNET_FLAG_TRANSFER_ASCII FTP_TRANSFER_TYPE_ASCII
#define FTP_TRANSFER_TYPE_BINARY 0x00000002
#define INTERNET_FLAG_TRANSFER_BINARY FTP_TRANSFER_TYPE_BINARY
#define _SECURITY_INTERNET_MASK INTERNET_FLAG_IGNORE_CERT_CN_INVALID | INTERNET_FLAG_IGNORE_CERT_DATE_INVALID | INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTPS | INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTP
#define _INTERNET_FLAGS_MASK INTERNET_FLAG_RELOAD | INTERNET_FLAG_RAW_DATA | INTERNET_FLAG_EXISTING_CONNECT | INTERNET_FLAG_ASYNC | INTERNET_FLAG_PASSIVE | INTERNET_FLAG_NO_CACHE_WRITE | INTERNET_FLAG_MAKE_PERSISTENT | INTERNET_FLAG_FROM_CACHE | INTERNET_FLAG_SECURE | INTERNET_FLAG_KEEP_CONNECTION | INTERNET_FLAG_NO_AUTO_REDIRECT | INTERNET_FLAG_READ_PREFETCH | INTERNET_FLAG_NO_COOKIES | INTERNET_FLAG_NO_AUTH | INTERNET_FLAG_CACHE_IF_NET_FAIL | _SECURITY_INTERNET_MASK | INTERNET_FLAG_RESYNCHRONIZE | INTERNET_FLAG_HYPERLINK | INTERNET_FLAG_NO_UI | INTERNET_FLAG_PRAGMA_NOCACHE | INTERNET_FLAG_CACHE_ASYNC | INTERNET_FLAG_FORMS_SUBMIT | INTERNET_FLAG_NEED_FILE | INTERNET_FLAG_RESTRICTED_ZONE | INTERNET_FLAG_TRANSFER_BINARY | INTERNET_FLAG_TRANSFER_ASCII | INTERNET_FLAG_FWD_BACK | INTERNET_FLAG_BGUPDATE
#define INTERNET_ERROR_MASK_INSERT_CDROM 0x1
#define INTERNET_ERROR_MASK_COMBINED_SEC_CERT 0x2
#define INTERNET_ERROR_MASK_NEED_MSN_SSPI_PKG 0X4
#define INTERNET_ERROR_MASK_LOGIN_FAILURE_DISPLAY_ENTITY_BODY 0x8
#define INTERNET_OPTIONS_MASK _NOT(_INTERNET_FLAGS_MASK)
#define WININET_API_FLAG_ASYNC 0x00000001
#define WININET_API_FLAG_SYNC 0x00000004
#define WININET_API_FLAG_USE_CONTEXT 0x00000008
#define INTERNET_NO_CALLBACK 0
#define INTERNET_SCHEME_PARTIAL -2
#define INTERNET_SCHEME_UNKNOWN -1
#define INTERNET_SCHEME_DEFAULT 0
#define INTERNET_SCHEME_FTP 1
#define INTERNET_SCHEME_GOPHER 2
#define INTERNET_SCHEME_HTTP 3
#define INTERNET_SCHEME_HTTPS 4
#define INTERNET_SCHEME_FILE 5
#define INTERNET_SCHEME_NEWS 6
#define INTERNET_SCHEME_MAILTO 7
#define INTERNET_SCHEME_SOCKS 8
#define INTERNET_SCHEME_JAVASCRIPT 9
#define INTERNET_SCHEME_VBSCRIPT 10
#define INTERNET_SCHEME_RES 11
#define INTERNET_SCHEME_FIRST INTERNET_SCHEME_FTP
#define INTERNET_SCHEME_LAST INTERNET_SCHEME_RES
#define INTERNET_PREFETCH_PROGRESS 0
#define INTERNET_PREFETCH_COMPLETE 1
#define INTERNET_PREFETCH_ABORTED 2
#define IDSI_FLAG_KEEP_ALIVE 0x00000001
#define IDSI_FLAG_SECURE 0x00000002
#define IDSI_FLAG_PROXY 0x00000004
#define IDSI_FLAG_TUNNEL 0x00000008
#define ISO_FORCE_DISCONNECTED 0x01
#define INTERNET_OPEN_TYPE_PRECONFIG 0
#define INTERNET_OPEN_TYPE_DIRECT 1
#define INTERNET_OPEN_TYPE_PROXY 3
#define INTERNET_OPEN_TYPE_PRECONFIG_WITH_NO_AUTOPROXY 4
#define PRE_CONFIG_INTERNET_ACCESS INTERNET_OPEN_TYPE_PRECONFIG
#define LOCAL_INTERNET_ACCESS INTERNET_OPEN_TYPE_DIRECT
#define GATEWAY_INTERNET_ACCESS 2
#define CERN_PROXY_INTERNET_ACCESS INTERNET_OPEN_TYPE_PROXY
#define INTERNET_SERVICE_FTP 1
#define INTERNET_SERVICE_GOPHER 2
#define INTERNET_SERVICE_HTTP 3
#define INTERNET_OPTION_CALLBACK 1
#define INTERNET_OPTION_CONNECT_TIMEOUT 2
#define INTERNET_OPTION_CONNECT_RETRIES 3
#define INTERNET_OPTION_CONNECT_BACKOFF 4
#define INTERNET_OPTION_SEND_TIMEOUT 5
#define INTERNET_OPTION_CONTROL_SEND_TIMEOUT INTERNET_OPTION_SEND_TIMEOUT
#define INTERNET_OPTION_RECEIVE_TIMEOUT 6
#define INTERNET_OPTION_CONTROL_RECEIVE_TIMEOUT INTERNET_OPTION_RECEIVE_TIMEOUT
#define INTERNET_OPTION_DATA_SEND_TIMEOUT 7
#define INTERNET_OPTION_DATA_RECEIVE_TIMEOUT 8
#define INTERNET_OPTION_HANDLE_TYPE 9
#define INTERNET_OPTION_LISTEN_TIMEOUT 11
#define INTERNET_OPTION_READ_BUFFER_SIZE 12
#define INTERNET_OPTION_WRITE_BUFFER_SIZE 13
#define INTERNET_OPTION_ASYNC_ID 15
#define INTERNET_OPTION_ASYNC_PRIORITY 16
#define INTERNET_OPTION_PARENT_HANDLE 21
#define INTERNET_OPTION_KEEP_CONNECTION 22
#define INTERNET_OPTION_REQUEST_FLAGS 23
#define INTERNET_OPTION_EXTENDED_ERROR 24
#define INTERNET_OPTION_OFFLINE_MODE 26
#define INTERNET_OPTION_CACHE_STREAM_HANDLE 27
#define INTERNET_OPTION_USERNAME 28
#define INTERNET_OPTION_PASSWORD 29
#define INTERNET_OPTION_ASYNC 30
#define INTERNET_OPTION_SECURITY_FLAGS 31
#define INTERNET_OPTION_SECURITY_CERTIFICATE_STRUCT 32
#define INTERNET_OPTION_DATAFILE_NAME 33
#define INTERNET_OPTION_URL 34
#define INTERNET_OPTION_SECURITY_CERTIFICATE 35
#define INTERNET_OPTION_SECURITY_KEY_BITNESS 36
#define INTERNET_OPTION_REFRESH 37
#define INTERNET_OPTION_PROXY 38
#define INTERNET_OPTION_SETTINGS_CHANGED 39
#define INTERNET_OPTION_VERSION 40
#define INTERNET_OPTION_USER_AGENT 41
#define INTERNET_OPTION_END_BROWSER_SESSION 42
#define INTERNET_OPTION_PROXY_USERNAME 43
#define INTERNET_OPTION_PROXY_PASSWORD 44
#define INTERNET_OPTION_CONTEXT_VALUE 45
#define INTERNET_OPTION_CONNECT_LIMIT 46
#define INTERNET_OPTION_SECURITY_SELECT_CLIENT_CERT 47
#define INTERNET_OPTION_POLICY 48
#define INTERNET_OPTION_DISCONNECTED_TIMEOUT 49
#define INTERNET_OPTION_CONNECTED_STATE 50
#define INTERNET_OPTION_IDLE_STATE 51
#define INTERNET_OPTION_OFFLINE_SEMANTICS 52
#define INTERNET_OPTION_SECONDARY_CACHE_KEY 53
#define INTERNET_OPTION_CALLBACK_FILTER 54
#define INTERNET_OPTION_CONNECT_TIME 55
#define INTERNET_OPTION_SEND_THROUGHPUT 56
#define INTERNET_OPTION_RECEIVE_THROUGHPUT 57
#define INTERNET_OPTION_REQUEST_PRIORITY 58
#define INTERNET_OPTION_HTTP_VERSION 59
#define INTERNET_OPTION_RESET_URLCACHE_SESSION 60
#define INTERNET_OPTION_ERROR_MASK 62
#define INTERNET_OPTION_FROM_CACHE_TIMEOUT 63
#define INTERNET_OPTION_BYPASS_EDITED_ENTRY 64
#define INTERNET_OPTION_DIAGNOSTIC_SOCKET_INFO 67
#define INTERNET_OPTION_CODEPAGE 68
#define INTERNET_OPTION_CACHE_TIMESTAMPS 69
#define INTERNET_OPTION_DISABLE_AUTODIAL 70
#define INTERNET_OPTION_MAX_CONNS_PER_SERVER 73
#define INTERNET_OPTION_MAX_CONNS_PER_1_0_SERVER 74
#define INTERNET_OPTION_PER_CONNECTION_OPTION 75
#define INTERNET_OPTION_DIGEST_AUTH_UNLOAD 76
#define INTERNET_OPTION_IGNORE_OFFLINE 77
#define INTERNET_OPTION_IDENTITY 78
#define INTERNET_OPTION_REMOVE_IDENTITY 79
#define INTERNET_OPTION_ALTER_IDENTITY 80
#define INTERNET_OPTION_SUPPRESS_BEHAVIOR 81
#define INTERNET_OPTION_AUTODIAL_MODE 82
#define INTERNET_OPTION_AUTODIAL_CONNECTION 83
#define INTERNET_OPTION_CLIENT_CERT_CONTEXT 84
#define INTERNET_OPTION_AUTH_FLAGS 85
#define INTERNET_OPTION_COOKIES_3RD_PARTY 86
#define INTERNET_OPTION_DISABLE_PASSPORT_AUTH 87
#define INTERNET_OPTION_SEND_UTF8_SERVERNAME_TO_PROXY 88
#define INTERNET_OPTION_EXEMPT_CONNECTION_LIMIT 89
#define INTERNET_OPTION_ENABLE_PASSPORT_AUTH 90
#define INTERNET_OPTION_HIBERNATE_INACTIVE_WORKER_THREADS 91
#define INTERNET_OPTION_ACTIVATE_WORKER_THREADS 92
#define INTERNET_OPTION_RESTORE_WORKER_THREAD_DEFAULTS 93
#define INTERNET_OPTION_SOCKET_SEND_BUFFER_LENGTH 94
#define INTERNET_OPTION_PROXY_SETTINGS_CHANGED 95
#define INTERNET_OPTION_DATAFILE_EXT 96
#define INTERNET_FIRST_OPTION INTERNET_OPTION_CALLBACK
#define INTERNET_LAST_OPTION INTERNET_OPTION_DATAFILE_EXT
#define INTERNET_PRIORITY_FOREGROUND 1000
#define INTERNET_HANDLE_TYPE_INTERNET 1
#define INTERNET_HANDLE_TYPE_CONNECT_FTP 2
#define INTERNET_HANDLE_TYPE_CONNECT_GOPHER 3
#define INTERNET_HANDLE_TYPE_CONNECT_HTTP 4
#define INTERNET_HANDLE_TYPE_FTP_FIND 5
#define INTERNET_HANDLE_TYPE_FTP_FIND_HTML 6
#define INTERNET_HANDLE_TYPE_FTP_FILE 7
#define INTERNET_HANDLE_TYPE_FTP_FILE_HTML 8
#define INTERNET_HANDLE_TYPE_GOPHER_FIND 9
#define INTERNET_HANDLE_TYPE_GOPHER_FIND_HTML 10
#define INTERNET_HANDLE_TYPE_GOPHER_FILE 11
#define INTERNET_HANDLE_TYPE_GOPHER_FILE_HTML 12
#define INTERNET_HANDLE_TYPE_HTTP_REQUEST 13
#define INTERNET_HANDLE_TYPE_FILE_REQUEST 14
#define AUTH_FLAG_DISABLE_NEGOTIATE 0x00000001
#define AUTH_FLAG_ENABLE_NEGOTIATE 0x00000002
#define AUTH_FLAG_DISABLE_BASIC_CLEARCHANNEL 0x00000004
#define SECURITY_FLAG_SECURE 0x00000001
#define SECURITY_FLAG_STRENGTH_WEAK 0x10000000
#define SECURITY_FLAG_STRENGTH_MEDIUM 0x40000000
#define SECURITY_FLAG_STRENGTH_STRONG 0x20000000
#define SECURITY_FLAG_UNKNOWNBIT 0x80000000
#define SECURITY_FLAG_FORTEZZA 0x08000000
#define SECURITY_FLAG_NORMALBITNESS SECURITY_FLAG_STRENGTH_WEAK
#define SECURITY_FLAG_SSL 0x00000002
#define SECURITY_FLAG_SSL3 0x00000004
#define SECURITY_FLAG_PCT 0x00000008
#define SECURITY_FLAG_PCT4 0x00000010
#define SECURITY_FLAG_IETFSSL4 0x00000020
#define SECURITY_FLAG_40BIT SECURITY_FLAG_STRENGTH_WEAK
#define SECURITY_FLAG_128BIT SECURITY_FLAG_STRENGTH_STRONG
#define SECURITY_FLAG_56BIT SECURITY_FLAG_STRENGTH_MEDIUM
#define SECURITY_FLAG_IGNORE_REVOCATION 0x00000080
#define SECURITY_FLAG_IGNORE_UNKNOWN_CA 0x00000100
#define SECURITY_FLAG_IGNORE_WRONG_USAGE 0x00000200
#define SECURITY_FLAG_IGNORE_CERT_CN_INVALID INTERNET_FLAG_IGNORE_CERT_CN_INVALID
#define SECURITY_FLAG_IGNORE_CERT_DATE_INVALID INTERNET_FLAG_IGNORE_CERT_DATE_INVALID
#define SECURITY_FLAG_IGNORE_REDIRECT_TO_HTTPS INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTPS
#define SECURITY_FLAG_IGNORE_REDIRECT_TO_HTTP INTERNET_FLAG_IGNORE_REDIRECT_TO_HTTP
#define AUTODIAL_MODE_NEVER 1
#define AUTODIAL_MODE_ALWAYS 2
#define AUTODIAL_MODE_NO_NETWORK_PRESENT 4
#define INTERNET_STATUS_RESOLVING_NAME 10
#define INTERNET_STATUS_NAME_RESOLVED 11
#define INTERNET_STATUS_CONNECTING_TO_SERVER 20
#define INTERNET_STATUS_CONNECTED_TO_SERVER 21
#define INTERNET_STATUS_SENDING_REQUEST 30
#define INTERNET_STATUS_REQUEST_SENT 31
#define INTERNET_STATUS_RECEIVING_RESPONSE 40
#define INTERNET_STATUS_RESPONSE_RECEIVED 41
#define INTERNET_STATUS_CTL_RESPONSE_RECEIVED 42
#define INTERNET_STATUS_PREFETCH 43
#define INTERNET_STATUS_CLOSING_CONNECTION 50
#define INTERNET_STATUS_CONNECTION_CLOSED 51
#define INTERNET_STATUS_HANDLE_CREATED 60
#define INTERNET_STATUS_HANDLE_CLOSING 70
#define INTERNET_STATUS_DETECTING_PROXY 80
#define INTERNET_STATUS_REQUEST_COMPLETE 100
#define INTERNET_STATUS_REDIRECT 110
#define INTERNET_STATUS_INTERMEDIATE_RESPONSE 120
#define INTERNET_STATUS_USER_INPUT_REQUIRED 140
#define INTERNET_STATUS_STATE_CHANGE 200
#define INTERNET_STATUS_COOKIE_SENT 320
#define INTERNET_STATUS_COOKIE_RECEIVED 321
#define INTERNET_STATUS_PRIVACY_IMPACTED 324
#define INTERNET_STATUS_P3P_HEADER 325
#define INTERNET_STATUS_P3P_POLICYREF 326
#define INTERNET_STATUS_COOKIE_HISTORY 327
#define INTERNET_STATE_CONNECTED 0x00000001
#define INTERNET_STATE_DISCONNECTED 0x00000002
#define INTERNET_STATE_DISCONNECTED_BY_USER 0x00000010
#define INTERNET_STATE_IDLE 0x00000100
#define INTERNET_STATE_BUSY 0x00000200
#define COOKIE_STATE_UNKNOWN 0x0
#define COOKIE_STATE_ACCEPT 0x1
#define COOKIE_STATE_PROMPT 0x2
#define COOKIE_STATE_LEASH 0x3
#define COOKIE_STATE_DOWNGRADE 0x4
#define COOKIE_STATE_REJECT 0x5
#define COOKIE_STATE_MAX COOKIE_STATE_REJECT
#define FTP_TRANSFER_TYPE_UNKNOWN 0x00000000
#define _FTP_TRANSFER_TYPE_MASK (FTP_TRANSFER_TYPE_ASCII | FTP_TRANSFER_TYPE_BINARY)
#define HTTP_MAJOR_VERSION 1
#define HTTP_MINOR_VERSION 0
#define HTTP_VERSION "HTTP/1.0"
#define HTTP_QUERY_MIME_VERSION 0
#define HTTP_QUERY_CONTENT_TYPE 1
#define HTTP_QUERY_CONTENT_TRANSFER_ENCODING 2
#define HTTP_QUERY_CONTENT_ID 3
#define HTTP_QUERY_CONTENT_DESCRIPTION 4
#define HTTP_QUERY_CONTENT_LENGTH 5
#define HTTP_QUERY_CONTENT_LANGUAGE 6
#define HTTP_QUERY_ALLOW 7
#define HTTP_QUERY_PUBLIC 8
#define HTTP_QUERY_DATE 9
#define HTTP_QUERY_EXPIRES 10
#define HTTP_QUERY_LAST_MODIFIED 11
#define HTTP_QUERY_MESSAGE_ID 12
#define HTTP_QUERY_URI 13
#define HTTP_QUERY_DERIVED_FROM 14
#define HTTP_QUERY_COST 15
#define HTTP_QUERY_LINK 16
#define HTTP_QUERY_PRAGMA 17
#define HTTP_QUERY_VERSION 18
#define HTTP_QUERY_STATUS_CODE 19
#define HTTP_QUERY_STATUS_TEXT 20
#define HTTP_QUERY_RAW_HEADERS 21
#define HTTP_QUERY_RAW_HEADERS_CRLF 22
#define HTTP_QUERY_CONNECTION 23
#define HTTP_QUERY_ACCEPT 24
#define HTTP_QUERY_ACCEPT_CHARSET 25
#define HTTP_QUERY_ACCEPT_ENCODING 26
#define HTTP_QUERY_ACCEPT_LANGUAGE 27
#define HTTP_QUERY_AUTHORIZATION 28
#define HTTP_QUERY_CONTENT_ENCODING 29
#define HTTP_QUERY_FORWARDED 30
#define HTTP_QUERY_FROM 31
#define HTTP_QUERY_IF_MODIFIED_SINCE 32
#define HTTP_QUERY_LOCATION 33
#define HTTP_QUERY_ORIG_URI 34
#define HTTP_QUERY_REFERER 35
#define HTTP_QUERY_RETRY_AFTER 36
#define HTTP_QUERY_SERVER 37
#define HTTP_QUERY_TITLE 38
#define HTTP_QUERY_USER_AGENT 39
#define HTTP_QUERY_WWW_AUTHENTICATE 40
#define HTTP_QUERY_PROXY_AUTHENTICATE 41
#define HTTP_QUERY_ACCEPT_RANGES 42
#define HTTP_QUERY_SET_COOKIE 43
#define HTTP_QUERY_COOKIE 44
#define HTTP_QUERY_REQUEST_METHOD 45
#define HTTP_QUERY_REFRESH 46
#define HTTP_QUERY_CONTENT_DISPOSITION 47
#define HTTP_QUERY_AGE 48
#define HTTP_QUERY_CACHE_CONTROL 49
#define HTTP_QUERY_CONTENT_BASE 50
#define HTTP_QUERY_CONTENT_LOCATION 51
#define HTTP_QUERY_CONTENT_MD5 52
#define HTTP_QUERY_CONTENT_RANGE 53
#define HTTP_QUERY_HOST 55
#define HTTP_QUERY_IF_MATCH 56
#define HTTP_QUERY_IF_NONE_MATCH 57
#define HTTP_QUERY_IF_RANGE 58
#define HTTP_QUERY_IF_UNMODIFIED_SINCE 59
#define HTTP_QUERY_MAX_FORWARDS 60
#define HTTP_QUERY_PROXY_AUTHORIZATION 61
#define HTTP_QUERY_RANGE 62
#define HTTP_QUERY_TRANSFER_ENCODING 63
#define HTTP_QUERY_UPGRADE 64
#define HTTP_QUERY_VARY 65
#define HTTP_QUERY_VIA 66
#define HTTP_QUERY_WARNING 67
#define HTTP_QUERY_EXPECT 68
#define HTTP_QUERY_PROXY_CONNECTION 69
#define HTTP_QUERY_UNLESS_MODIFIED_SINCE 70
#define HTTP_QUERY_ECHO_REQUEST 71
#define HTTP_QUERY_ECHO_REPLY 72
#define HTTP_QUERY_ECHO_HEADERS 73
#define HTTP_QUERY_ECHO_HEADERS_CRLF 74
#define HTTP_QUERY_PROXY_SUPPORT 75
#define HTTP_QUERY_AUTHENTICATION_INFO 76
#define HTTP_QUERY_PASSPORT_URLS 77
#define HTTP_QUERY_PASSPORT_CONFIG 78
#define HTTP_QUERY_CUSTOM 65535
#define HTTP_QUERY_FLAG_REQUEST_HEADERS 0x80000000
#define HTTP_QUERY_FLAG_SYSTEMTIME 0x40000000
#define HTTP_QUERY_FLAG_NUMBER 0x20000000
#define HTTP_QUERY_FLAG_COALESCE 0x10000000
#define HTTP_QUERY_MODIFIER_FLAGS_MASK (HTTP_QUERY_FLAG_REQUEST_HEADERS | HTTP_QUERY_FLAG_SYSTEMTIME | HTTP_QUERY_FLAG_NUMBER | HTTP_QUERY_FLAG_COALESCE )
#define HTTP_STATUS_CONTINUE 100
#define HTTP_STATUS_SWITCH_PROTOCOLS 101
#define HTTP_STATUS_OK 200
#define HTTP_STATUS_CREATED 201
#define HTTP_STATUS_ACCEPTED 202
#define HTTP_STATUS_PARTIAL 203
#define HTTP_STATUS_NO_CONTENT 204
#define HTTP_STATUS_RESET_CONTENT 205
#define HTTP_STATUS_PARTIAL_CONTENT 206
#define HTTP_STATUS_AMBIGUOUS 300
#define HTTP_STATUS_MOVED 301
#define HTTP_STATUS_REDIRECT 302
#define HTTP_STATUS_REDIRECT_METHOD 303
#define HTTP_STATUS_NOT_MODIFIED 304
#define HTTP_STATUS_USE_PROXY 305
#define HTTP_STATUS_REDIRECT_KEEP_VERB 307
#define HTTP_STATUS_BAD_REQUEST 400
#define HTTP_STATUS_DENIED 401
#define HTTP_STATUS_PAYMENT_REQ 402
#define HTTP_STATUS_FORBIDDEN 403
#define HTTP_STATUS_NOT_FOUND 404
#define HTTP_STATUS_BAD_METHOD 405
#define HTTP_STATUS_NONE_ACCEPTABLE 406
#define HTTP_STATUS_PROXY_AUTH_REQ 407
#define HTTP_STATUS_REQUEST_TIMEOUT 408
#define HTTP_STATUS_CONFLICT 409
#define HTTP_STATUS_GONE 410
#define HTTP_STATUS_AUTH_REFUSED 411
#define HTTP_STATUS_PRECOND_FAILED 412
#define HTTP_STATUS_REQUEST_TOO_LARGE 413
#define HTTP_STATUS_URI_TOO_LONG 414
#define HTTP_STATUS_UNSUPPORTED_MEDIA 415
#define HTTP_STATUS_RETRY_WITH 449
#define HTTP_STATUS_SERVER_ERROR 500
#define HTTP_STATUS_NOT_SUPPORTED 501
#define HTTP_STATUS_BAD_GATEWAY 502
#define HTTP_STATUS_SERVICE_UNAVAIL 503
#define HTTP_STATUS_GATEWAY_TIMEOUT 504
#define HTTP_STATUS_VERSION_NOT_SUP 505
#define HTTP_STATUS_FIRST HTTP_STATUS_CONTINUE
#define HTTP_STATUS_LAST HTTP_STATUS_VERSION_NOT_SUP
#define HTTP_ADDREQ_INDEX_MASK 0x0000FFFF
#define HTTP_ADDREQ_FLAGS_MASK 0xFFFF0000
#define HTTP_ADDREQ_FLAG_ADD_IF_NEW 0x10000000
#define HTTP_ADDREQ_FLAG_ADD 0x20000000
#define HTTP_ADDREQ_FLAG_COALESCE_WITH_COMMA 0x40000000
#define HTTP_ADDREQ_FLAG_COALESCE_WITH_SEMICOLON 0x01000000
#define HTTP_ADDREQ_FLAG_COALESCE HTTP_ADDREQ_FLAG_COALESCE_WITH_COMMA
#define HTTP_ADDREQ_FLAG_REPLACE 0x80000000
#define HSR_ASYNC WININET_API_FLAG_ASYNC
#define HSR_SYNC WININET_API_FLAG_SYNC
#define HSR_USE_CONTEXT WININET_API_FLAG_USE_CONTEXT
#define HSR_INITIATE 0x00000008
#define HSR_DOWNLOAD 0x00000010
#define HSR_CHUNKED 0x00000020
#define INTERNET_ERROR_BASE 12000
#define ERROR_INTERNET_OUT_OF_HANDLES (INTERNET_ERROR_BASE + 1)
#define ERROR_INTERNET_TIMEOUT (INTERNET_ERROR_BASE + 2)
#define ERROR_INTERNET_EXTENDED_ERROR (INTERNET_ERROR_BASE + 3)
#define ERROR_INTERNET_INTERNAL_ERROR (INTERNET_ERROR_BASE + 4)
#define ERROR_INTERNET_INVALID_URL (INTERNET_ERROR_BASE + 5)
#define ERROR_INTERNET_UNRECOGNIZED_SCHEME (INTERNET_ERROR_BASE + 6)
#define ERROR_INTERNET_NAME_NOT_RESOLVED (INTERNET_ERROR_BASE + 7)
#define ERROR_INTERNET_PROTOCOL_NOT_FOUND (INTERNET_ERROR_BASE + 8)
#define ERROR_INTERNET_INVALID_OPTION (INTERNET_ERROR_BASE + 9)
#define ERROR_INTERNET_BAD_OPTION_LENGTH (INTERNET_ERROR_BASE + 10)
#define ERROR_INTERNET_OPTION_NOT_SETTABLE (INTERNET_ERROR_BASE + 11)
#define ERROR_INTERNET_SHUTDOWN (INTERNET_ERROR_BASE + 12)
#define ERROR_INTERNET_INCORRECT_USER_NAME (INTERNET_ERROR_BASE + 13)
#define ERROR_INTERNET_INCORRECT_PASSWORD (INTERNET_ERROR_BASE + 14)
#define ERROR_INTERNET_LOGIN_FAILURE (INTERNET_ERROR_BASE + 15)
#define ERROR_INTERNET_INVALID_OPERATION (INTERNET_ERROR_BASE + 16)
#define ERROR_INTERNET_OPERATION_CANCELLED (INTERNET_ERROR_BASE + 17)
#define ERROR_INTERNET_INCORRECT_HANDLE_TYPE (INTERNET_ERROR_BASE + 18)
#define ERROR_INTERNET_INCORRECT_HANDLE_STATE (INTERNET_ERROR_BASE + 19)
#define ERROR_INTERNET_NOT_PROXY_REQUEST (INTERNET_ERROR_BASE + 20)
#define ERROR_INTERNET_REGISTRY_VALUE_NOT_FOUND (INTERNET_ERROR_BASE + 21)
#define ERROR_INTERNET_BAD_REGISTRY_PARAMETER (INTERNET_ERROR_BASE + 22)
#define ERROR_INTERNET_NO_DIRECT_ACCESS (INTERNET_ERROR_BASE + 23)
#define ERROR_INTERNET_NO_CONTEXT (INTERNET_ERROR_BASE + 24)
#define ERROR_INTERNET_NO_CALLBACK (INTERNET_ERROR_BASE + 25)
#define ERROR_INTERNET_REQUEST_PENDING (INTERNET_ERROR_BASE + 26)
#define ERROR_INTERNET_INCORRECT_FORMAT (INTERNET_ERROR_BASE + 27)
#define ERROR_INTERNET_ITEM_NOT_FOUND (INTERNET_ERROR_BASE + 28)
#define ERROR_INTERNET_CANNOT_CONNECT (INTERNET_ERROR_BASE + 29)
#define ERROR_INTERNET_CONNECTION_ABORTED (INTERNET_ERROR_BASE + 30)
#define ERROR_INTERNET_CONNECTION_RESET (INTERNET_ERROR_BASE + 31)
#define ERROR_INTERNET_FORCE_RETRY (INTERNET_ERROR_BASE + 32)
#define ERROR_INTERNET_INVALID_PROXY_REQUEST (INTERNET_ERROR_BASE + 33)
#define ERROR_INTERNET_NEED_UI (INTERNET_ERROR_BASE + 34)
#define ERROR_INTERNET_HANDLE_EXISTS (INTERNET_ERROR_BASE + 36)
#define ERROR_INTERNET_SEC_CERT_DATE_INVALID (INTERNET_ERROR_BASE + 37)
#define ERROR_INTERNET_SEC_CERT_CN_INVALID (INTERNET_ERROR_BASE + 38)
#define ERROR_INTERNET_HTTP_TO_HTTPS_ON_REDIR (INTERNET_ERROR_BASE + 39)
#define ERROR_INTERNET_HTTPS_TO_HTTP_ON_REDIR (INTERNET_ERROR_BASE + 40)
#define ERROR_INTERNET_MIXED_SECURITY (INTERNET_ERROR_BASE + 41)
#define ERROR_INTERNET_CHG_POST_IS_NON_SECURE (INTERNET_ERROR_BASE + 42)
#define ERROR_INTERNET_POST_IS_NON_SECURE (INTERNET_ERROR_BASE + 43)
#define ERROR_INTERNET_CLIENT_AUTH_CERT_NEEDED (INTERNET_ERROR_BASE + 44)
#define ERROR_INTERNET_INVALID_CA (INTERNET_ERROR_BASE + 45)
#define ERROR_INTERNET_CLIENT_AUTH_NOT_SETUP (INTERNET_ERROR_BASE + 46)
#define ERROR_INTERNET_ASYNC_THREAD_FAILED (INTERNET_ERROR_BASE + 47)
#define ERROR_INTERNET_REDIRECT_SCHEME_CHANGE (INTERNET_ERROR_BASE + 48)
#define ERROR_INTERNET_DIALOG_PENDING (INTERNET_ERROR_BASE + 49)
#define ERROR_INTERNET_RETRY_DIALOG ( INTERNET_ERROR_BASE + 50)
#define ERROR_INTERNET_HTTPS_HTTP_SUBMIT_REDIR (INTERNET_ERROR_BASE + 52)
#define ERROR_INTERNET_INSERT_CDROM (INTERNET_ERROR_BASE + 53)
#define ERROR_INTERNET_FORTEZZA_LOGIN_NEEDED (INTERNET_ERROR_BASE + 54)
#define ERROR_INTERNET_SEC_CERT_ERRORS (INTERNET_ERROR_BASE + 55)
#define ERROR_INTERNET_SEC_CERT_NO_REV (INTERNET_ERROR_BASE + 56)
#define ERROR_INTERNET_SEC_CERT_REV_FAILED (INTERNET_ERROR_BASE + 57)
#define ERROR_FTP_TRANSFER_IN_PROGRESS (INTERNET_ERROR_BASE + 110)
#define ERROR_FTP_DROPPED (INTERNET_ERROR_BASE + 111)
#define ERROR_FTP_NO_PASSIVE_MODE (INTERNET_ERROR_BASE + 112)
#define ERROR_GOPHER_PROTOCOL_ERROR (INTERNET_ERROR_BASE + 130)
#define ERROR_GOPHER_NOT_FILE (INTERNET_ERROR_BASE + 131)
#define ERROR_GOPHER_DATA_ERROR (INTERNET_ERROR_BASE + 132)
#define ERROR_GOPHER_END_OF_DATA (INTERNET_ERROR_BASE + 133)
#define ERROR_GOPHER_INVALID_LOCATOR (INTERNET_ERROR_BASE + 134)
#define ERROR_GOPHER_INCORRECT_LOCATOR_TYPE (INTERNET_ERROR_BASE + 135)
#define ERROR_GOPHER_NOT_GOPHER_PLUS (INTERNET_ERROR_BASE + 136)
#define ERROR_GOPHER_ATTRIBUTE_NOT_FOUND (INTERNET_ERROR_BASE + 137)
#define ERROR_GOPHER_UNKNOWN_LOCATOR (INTERNET_ERROR_BASE + 138)
#define ERROR_HTTP_HEADER_NOT_FOUND (INTERNET_ERROR_BASE + 150)
#define ERROR_HTTP_DOWNLEVEL_SERVER (INTERNET_ERROR_BASE + 151)
#define ERROR_HTTP_INVALID_SERVER_RESPONSE (INTERNET_ERROR_BASE + 152)
#define ERROR_HTTP_INVALID_HEADER (INTERNET_ERROR_BASE + 153)
#define ERROR_HTTP_INVALID_QUERY_REQUEST (INTERNET_ERROR_BASE + 154)
#define ERROR_HTTP_HEADER_ALREADY_EXISTS (INTERNET_ERROR_BASE + 155)
#define ERROR_HTTP_REDIRECT_FAILED (INTERNET_ERROR_BASE + 156)
#define ERROR_HTTP_NOT_REDIRECTED (INTERNET_ERROR_BASE + 160)
#define ERROR_HTTP_COOKIE_NEEDS_CONFIRMATION (INTERNET_ERROR_BASE + 161)
#define ERROR_HTTP_COOKIE_DECLINED (INTERNET_ERROR_BASE + 162)
#define ERROR_HTTP_REDIRECT_NEEDS_CONFIRMATION (INTERNET_ERROR_BASE + 168)
#define ERROR_INTERNET_SECURITY_CHANNEL_ERROR (INTERNET_ERROR_BASE + 157)
#define ERROR_INTERNET_UNABLE_TO_CACHE_FILE (INTERNET_ERROR_BASE + 158)
#define ERROR_INTERNET_TCPIP_NOT_INSTALLED (INTERNET_ERROR_BASE + 159)
#define ERROR_INTERNET_DISCONNECTED (INTERNET_ERROR_BASE + 163)
#define ERROR_INTERNET_SERVER_UNREACHABLE (INTERNET_ERROR_BASE + 164)
#define ERROR_INTERNET_PROXY_SERVER_UNREACHABLE (INTERNET_ERROR_BASE + 165)
#define ERROR_INTERNET_BAD_AUTO_PROXY_SCRIPT (INTERNET_ERROR_BASE + 166)
#define ERROR_INTERNET_UNABLE_TO_DOWNLOAD_SCRIPT (INTERNET_ERROR_BASE + 167)
#define ERROR_INTERNET_SEC_INVALID_CERT (INTERNET_ERROR_BASE + 169)
#define ERROR_INTERNET_SEC_CERT_REVOKED (INTERNET_ERROR_BASE + 170)
#define ERROR_INTERNET_FAILED_DUETOSECURITYCHECK (INTERNET_ERROR_BASE + 171)
#define ERROR_INTERNET_NOT_INITIALIZED (INTERNET_ERROR_BASE + 172)
#define ERROR_INTERNET_NEED_MSN_SSPI_PKG (INTERNET_ERROR_BASE + 173)
#define ERROR_INTERNET_LOGIN_FAILURE_DISPLAY_ENTITY_BODY (INTERNET_ERROR_BASE + 174)
#define INTERNET_ERROR_LAST ERROR_INTERNET_LOGIN_FAILURE_DISPLAY_ENTITY_BODY
#define FLAG_ICC_FORCE_CONNECTION 0x00000001
#define INTERNET_AUTODIAL_FORCE_ONLINE 1
#define INTERNET_AUTODIAL_FORCE_UNATTENDED 2
#define INTERNET_AUTODIAL_FAILIFSECURITYCHECK 4
#define INTERNET_AUTODIAL_OVERRIDE_NET_PRESENT 8
#define INTERNET_CONNECTION_MODEM 0x01
#define INTERNET_CONNECTION_LAN 0x02
#define INTERNET_CONNECTION_PROXY 0x04
#define INTERNET_CONNECTION_MODEM_BUSY 0x08 
#define INTERNET_RAS_INSTALLED 0x10
#define INTERNET_CONNECTION_OFFLINE 0x20
#define INTERNET_CONNECTION_CONFIGURED 0x40
#define INTERNET_CUSTOMDIAL_CONNECT 0
#define INTERNET_CUSTOMDIAL_UNATTENDED 1
#define INTERNET_CUSTOMDIAL_DISCONNECT 2
#define INTERNET_CUSTOMDIAL_SHOWOFFLINE 4
#define INTERNET_CUSTOMDIAL_SAFE_FOR_UNATTENDED 1
#define INTERNET_CUSTOMDIAL_WILL_SUPPLY_STATE 2
#define INTERNET_CUSTOMDIAL_CAN_HANGUP 4
#define INTERNET_IDENTITY_FLAG_PRIVATE_CACHE 0x01
#define INTERNET_IDENTITY_FLAG_SHARED_CACHE 0x02
#define INTERNET_IDENTITY_FLAG_CLEAR_DATA 0x04
#define INTERNET_IDENTITY_FLAG_CLEAR_COOKIES 0x08
#define INTERNET_IDENTITY_FLAG_CLEAR_HISTORY 0x10
#define INTERNET_IDENTITY_FLAG_CLEAR_CONTENT 0x20
#define INTERNET_SUPPRESS_RESET_ALL 0x00
#define INTERNET_SUPPRESS_COOKIE_POLICY 0x01
#define INTERNET_SUPPRESS_COOKIE_POLICY_RESET 0x02
#define PRIVACY_TEMPLATE_NO_COOKIES 0
#define PRIVACY_TEMPLATE_HIGH 1
#define PRIVACY_TEMPLATE_MEDIUM_HIGH 2
#define PRIVACY_TEMPLATE_MEDIUM 3
#define PRIVACY_TEMPLATE_MEDIUM_LOW 4
#define PRIVACY_TEMPLATE_LOW 5
#define PRIVACY_TEMPLATE_CUSTOM 100
#define PRIVACY_TEMPLATE_ADVANCED 101
#define PRIVACY_TEMPLATE_MAX PRIVACY_TEMPLATE_LOW
#define PRIVACY_TYPE_FIRST_PARTY 0
#define PRIVACY_TYPE_THIRD_PARTY 1
#define WNNC_NET_MSNET 0x00010000
#define WNNC_NET_LANMAN 0x00020000
#define WNNC_NET_NETWARE 0x00030000
#define WNNC_NET_VINES 0x00040000
#define WNNC_NET_10NET 0x00050000
#define WNNC_NET_LOCUS 0x00060000
#define WNNC_NET_SUN_PC_NFS 0x00070000
#define WNNC_NET_LANSTEP 0x00080000
#define WNNC_NET_9TILES 0x00090000
#define WNNC_NET_LANTASTIC 0x000A0000
#define WNNC_NET_AS400 0x000B0000
#define WNNC_NET_FTP_NFS 0x000C0000
#define WNNC_NET_PATHWORKS 0x000D0000
#define WNNC_NET_LIFENET 0x000E0000
#define WNNC_NET_POWERLAN 0x000F0000
#define WNNC_NET_BWNFS 0x00100000
#define WNNC_NET_COGENT 0x00110000
#define WNNC_NET_FARALLON 0x00120000
#define WNNC_NET_APPLETALK 0x00130000
#define RESOURCE_CONNECTED 0x00000001
#define RESOURCE_GLOBALNET 0x00000002
#define RESOURCE_REMEMBERED 0x00000003
#define RESOURCE_RECENT 0x00000004
#define RESOURCE_CONTEXT 0x00000005
#define RESOURCETYPE_ANY 0x00000000
#define RESOURCETYPE_DISK 0x00000001
#define RESOURCETYPE_PRINT 0x00000002
#define RESOURCETYPE_RESERVED 0x00000008
#define RESOURCETYPE_UNKNOWN 0xFFFFFFFF
#define RESOURCEUSAGE_CONNECTABLE 0x00000001
#define RESOURCEUSAGE_CONTAINER 0x00000002
#define RESOURCEUSAGE_NOLOCALDEVICE 0x00000004
#define RESOURCEUSAGE_SIBLING 0x00000008
#define RESOURCEUSAGE_ALL 0x00000003
#define RESOURCEUSAGE_RESERVED 0x80000000
#define RESOURCEDISPLAYTYPE_GENERIC 0x00000000
#define RESOURCEDISPLAYTYPE_DOMAIN 0x00000001
#define RESOURCEDISPLAYTYPE_SERVER 0x00000002
#define RESOURCEDISPLAYTYPE_SHARE 0x00000003
#define RESOURCEDISPLAYTYPE_FILE 0x00000004
#define RESOURCEDISPLAYTYPE_GROUP 0x00000005
#define RESOURCEDISPLAYTYPE_NETWORK 0x00000006
#define RESOURCEDISPLAYTYPE_ROOT 0x00000007
#define RESOURCEDISPLAYTYPE_SHAREADMIN 0x00000008
#define RESOURCEDISPLAYTYPE_DIRECTORY 0x00000009
#define RESOURCEDISPLAYTYPE_TREE 0x0000000A
#define NETPROPERTY_PERSISTENT 1
#define CONNECT_UPDATE_PROFILE 0x00000001
#define CONNECT_UPDATE_RECENT 0x00000002
#define CONNECT_TEMPORARY 0x00000004
#define CONNECT_INTERACTIVE 0x00000008
#define CONNECT_PROMPT 0x00000010
#define CONNECT_NEED_DRIVE 0x00000020
#define CONNECT_REFCOUNT 0x00000040
#define CONNECT_REDIRECT 0x00000080
#define CONNECT_LOCALDRIVE 0x00000100
#define CONNECT_CURRENT_MEDIA 0x00000200
#define CONNDLG_RO_PATH 0x00000001
#define CONNDLG_CONN_POINT 0x00000002
#define CONNDLG_USE_MRU 0x00000004
#define CONNDLG_HIDE_BOX 0x00000008
#define CONNDLG_PERSIST 0x00000010
#define CONNDLG_NOT_PERSIST 0x00000020
#define DISC_UPDATE_PROFILE 0x00000001
#define DISC_NO_FORCE 0x00000040
#define UNIVERSAL_NAME_INFO_LEVEL 0x00000001
#define REMOTE_NAME_INFO_LEVEL 0x00000002
#define WNFMT_MULTILINE 0x01
#define WNFMT_ABBREVIATED 0x02
#define WNFMT_INENUM 0x10
#define WNFMT_CONNECTION 0x20
#define NETINFO_DLL16 0x00000001
#define NETINFO_DISKRED 0x00000004
#define NETINFO_PRINTERRED 0x00000008
#define RP_LOGON 0x01
#define RP_INIFILE 0x02
#define PP_DISPLAYERRORS 0x01
#define WN_SUCCESS NO_ERROR
#define WN_NO_ERROR NO_ERROR
#define WN_NOT_SUPPORTED ERROR_NOT_SUPPORTED
#define WN_CANCEL ERROR_CANCELLED
#define WN_RETRY ERROR_RETRY
#define WN_NET_ERROR ERROR_UNEXP_NET_ERR
#define WN_MORE_DATA ERROR_MORE_DATA
#define WN_BAD_POINTER ERROR_INVALID_ADDRESS
#define WN_BAD_VALUE ERROR_INVALID_PARAMETER
#define WN_BAD_USER ERROR_BAD_USERNAME
#define WN_BAD_PASSWORD ERROR_INVALID_PASSWORD
#define WN_ACCESS_DENIED ERROR_ACCESS_DENIED
#define WN_FUNCTION_BUSY ERROR_BUSY
#define WN_WINDOWS_ERROR ERROR_UNEXP_NET_ERR
#define WN_OUT_OF_MEMORY ERROR_NOT_ENOUGH_MEMORY
#define WN_NO_NETWORK ERROR_NO_NETWORK
#define WN_EXTENDED_ERROR ERROR_EXTENDED_ERROR
#define WN_BAD_LEVEL ERROR_INVALID_LEVEL
#define WN_BAD_HANDLE ERROR_INVALID_HANDLE
#define WN_NOT_INITIALIZING ERROR_ALREADY_INITIALIZED
#define WN_NO_MORE_DEVICES ERROR_NO_MORE_DEVICES
#define WN_NOT_CONNECTED ERROR_NOT_CONNECTED
#define WN_OPEN_FILES ERROR_OPEN_FILES
#define WN_DEVICE_IN_USE ERROR_DEVICE_IN_USE
#define WN_BAD_NETNAME ERROR_BAD_NET_NAME
#define WN_BAD_LOCALNAME ERROR_BAD_DEVICE
#define WN_ALREADY_CONNECTED ERROR_ALREADY_ASSIGNED
#define WN_DEVICE_ERROR ERROR_GEN_FAILURE
#define WN_CONNECTION_CLOSED ERROR_CONNECTION_UNAVAIL
#define WN_NO_NET_OR_BAD_PATH ERROR_NO_NET_OR_BAD_PATH
#define WN_BAD_PROVIDER ERROR_BAD_PROVIDER
#define WN_CANNOT_OPEN_PROFILE ERROR_CANNOT_OPEN_PROFILE
#define WN_BAD_PROFILE ERROR_BAD_PROFILE
#define WN_BAD_DEV_TYPE ERROR_BAD_DEV_TYPE
#define WN_DEVICE_ALREADY_REMEMBERED ERROR_DEVICE_ALREADY_REMEMBERED
#define WN_NO_MORE_ENTRIES ERROR_NO_MORE_ITEMS
#define WN_NOT_CONTAINER ERROR_NOT_CONTAINER
#define WN_NOT_AUTHENTICATED ERROR_NOT_AUTHENTICATED
#define WN_NOT_LOGGED_ON ERROR_NOT_LOGGED_ON
#define WN_NOT_VALIDATED ERROR_NO_LOGON_SERVERS
#define WNCON_FORNETCARD 0x00000001
#define WNCON_NOTROUTED 0x00000002
#define WNCON_SLOWLINK 0x00000004
#define WNCON_DYNAMIC 0x00000008
#define MAX_LEADBYTES 12
#define MAX_DEFAULTCHAR 2
#define MB_PRECOMPOSED 0x00000001
#define MB_COMPOSITE 0x00000002
#define MB_USEGLYPHCHARS 0x00000004
#define MB_ERR_INVALID_CHARS 0x00000008
#define WC_DEFAULTCHECK 0x00000100
#define WC_COMPOSITECHECK 0x00000200
#define WC_DISCARDNS 0x00000010
#define WC_SEPCHARS 0x00000020
#define WC_DEFAULTCHAR 0x00000040
#define CT_CTYPE1 0x00000001
#define CT_CTYPE2 0x00000002
#define CT_CTYPE3 0x00000004
#define C1_UPPER 0x0001
#define C1_LOWER 0x0002
#define C1_DIGIT 0x0004
#define C1_SPACE 0x0008
#define C1_PUNCT 0x0010
#define C1_CNTRL 0x0020
#define C1_BLANK 0x0040
#define C1_XDIGIT 0x0080
#define C1_ALPHA 0x0100
#define C2_LEFTTORIGHT 0x0001
#define C2_RIGHTTOLEFT 0x0002
#define C2_EUROPENUMBER 0x0003
#define C2_EUROPESEPARATOR 0x0004
#define C2_EUROPETERMINATOR 0x0005
#define C2_ARABICNUMBER 0x0006
#define C2_COMMONSEPARATOR 0x0007
#define C2_BLOCKSEPARATOR 0x0008
#define C2_SEGMENTSEPARATOR 0x0009
#define C2_WHITESPACE 0x000A
#define C2_OTHERNEUTRAL 0x000B
#define C2_NOTAPPLICABLE 0x0000
#define C3_NONSPACING 0x0001
#define C3_DIACRITIC 0x0002
#define C3_VOWELMARK 0x0004
#define C3_SYMBOL 0x0008
#define C3_KATAKANA 0x0010
#define C3_HIRAGANA 0x0020
#define C3_HALFWIDTH 0x0040
#define C3_FULLWIDTH 0x0080
#define C3_IDEOGRAPH 0x0100
#define C3_KASHIDA 0x0200
#define C3_LEXICAL 0x0400
#define C3_ALPHA 0x8000
#define C3_NOTAPPLICABLE 0x0000
#define NORM_IGNORECASE 0x00000001
#define NORM_IGNORENONSPACE 0x00000002
#define NORM_IGNORESYMBOLS 0x00000004
#define NORM_IGNOREKANATYPE 0x00010000
#define NORM_IGNOREWIDTH 0x00020000
#define MAP_FOLDCZONE 0x00000010
#define MAP_PRECOMPOSED 0x00000020
#define MAP_COMPOSITE 0x00000040
#define MAP_FOLDDIGITS 0x00000080
#define LCMAP_LOWERCASE 0x00000100
#define LCMAP_UPPERCASE 0x00000200
#define LCMAP_SORTKEY 0x00000400
#define LCMAP_BYTEREV 0x00000800
#define LCMAP_HIRAGANA 0x00100000
#define LCMAP_KATAKANA 0x00200000
#define LCMAP_HALFWIDTH 0x00400000
#define LCMAP_FULLWIDTH 0x00800000
#define LCID_INSTALLED 0x00000001
#define LCID_SUPPORTED 0x00000002
#define CP_INSTALLED 0x00000001
#define CP_SUPPORTED 0x00000002
#define SORT_STRINGSORT 0x00001000
#define CP_ACP 0
#define CP_OEMCP 1
#define CP_MACCP 2
#define CTRY_DEFAULT 0
#define CTRY_AUSTRALIA 61
#define CTRY_AUSTRIA 43
#define CTRY_BELGIUM 32
#define CTRY_BRAZIL 55
#define CTRY_BULGARIA 359
#define CTRY_CANADA 2
#define CTRY_CROATIA 385
#define CTRY_CZECH 42
#define CTRY_DENMARK 45
#define CTRY_FINLAND 358
#define CTRY_FRANCE 33
#define CTRY_GERMANY 49
#define CTRY_GREECE 30
#define CTRY_HONG_KONG 852
#define CTRY_HUNGARY 36
#define CTRY_ICELAND 354
#define CTRY_IRELAND 353
#define CTRY_ITALY 39
#define CTRY_JAPAN 81
#define CTRY_MEXICO 52
#define CTRY_NETHERLANDS 31
#define CTRY_NEW_ZEALAND 64
#define CTRY_NORWAY 47
#define CTRY_POLAND 48
#define CTRY_PORTUGAL 351
#define CTRY_PRCHINA 86
#define CTRY_ROMANIA 40
#define CTRY_RUSSIA 7
#define CTRY_SINGAPORE 65
#define CTRY_SLOVAK 42
#define CTRY_SLOVENIA 386
#define CTRY_SOUTH_KOREA 82
#define CTRY_SPAIN 34
#define CTRY_SWEDEN 46
#define CTRY_SWITZERLAND 41
#define CTRY_TAIWAN 886
#define CTRY_TURKEY 90
#define CTRY_UNITED_KINGDOM 44
#define CTRY_UNITED_STATES 1
#define LOCALE_NOUSEROVERRIDE 0x80000000
#define LOCALE_USE_CP_ACP 0x40000000
#define LOCALE_ILANGUAGE 0x00000001
#define LOCALE_SLANGUAGE 0x00000002
#define LOCALE_SENGLANGUAGE 0x00001001
#define LOCALE_SABBREVLANGNAME 0x00000003
#define LOCALE_SNATIVELANGNAME 0x00000004
#define LOCALE_ICOUNTRY 0x00000005
#define LOCALE_SCOUNTRY 0x00000006
#define LOCALE_SENGCOUNTRY 0x00001002
#define LOCALE_SABBREVCTRYNAME 0x00000007
#define LOCALE_SNATIVECTRYNAME 0x00000008
#define LOCALE_IDEFAULTLANGUAGE 0x00000009
#define LOCALE_IDEFAULTCOUNTRY 0x0000000A
#define LOCALE_IDEFAULTCODEPAGE 0x0000000B
#define LOCALE_IDEFAULTANSICODEPAGE 0x00001004
#define LOCALE_SLIST 0x0000000C
#define LOCALE_IMEASURE 0x0000000D
#define LOCALE_SDECIMAL 0x0000000E
#define LOCALE_STHOUSAND 0x0000000F
#define LOCALE_SGROUPING 0x00000010
#define LOCALE_IDIGITS 0x00000011
#define LOCALE_ILZERO 0x00000012
#define LOCALE_INEGNUMBER 0x00001010
#define LOCALE_SNATIVEDIGITS 0x00000013
#define LOCALE_SCURRENCY 0x00000014
#define LOCALE_SINTLSYMBOL 0x00000015
#define LOCALE_SMONDECIMALSEP 0x00000016
#define LOCALE_SMONTHOUSANDSEP 0x00000017
#define LOCALE_SMONGROUPING 0x00000018
#define LOCALE_ICURRDIGITS 0x00000019
#define LOCALE_IINTLCURRDIGITS 0x0000001A
#define LOCALE_ICURRENCY 0x0000001B
#define LOCALE_INEGCURR 0x0000001C
#define LOCALE_SDATE 0x0000001D
#define LOCALE_STIME 0x0000001E
#define LOCALE_SSHORTDATE 0x0000001F
#define LOCALE_SLONGDATE 0x00000020
#define LOCALE_STIMEFORMAT 0x00001003
#define LOCALE_IDATE 0x00000021
#define LOCALE_ILDATE 0x00000022
#define LOCALE_ITIME 0x00000023
#define LOCALE_ITIMEMARKPOSN 0x00001005
#define LOCALE_ICENTURY 0x00000024
#define LOCALE_ITLZERO 0x00000025
#define LOCALE_IDAYLZERO 0x00000026
#define LOCALE_IMONLZERO 0x00000027
#define LOCALE_S1159 0x00000028
#define LOCALE_S2359 0x00000029
#define LOCALE_ICALENDARTYPE 0x00001009
#define LOCALE_IOPTIONALCALENDAR 0x0000100B
#define LOCALE_IFIRSTDAYOFWEEK 0x0000100C
#define LOCALE_IFIRSTWEEKOFYEAR 0x0000100D
#define LOCALE_SDAYNAME1 0x0000002A
#define LOCALE_SDAYNAME2 0x0000002B
#define LOCALE_SDAYNAME3 0x0000002C
#define LOCALE_SDAYNAME4 0x0000002D
#define LOCALE_SDAYNAME5 0x0000002E
#define LOCALE_SDAYNAME6 0x0000002F
#define LOCALE_SDAYNAME7 0x00000030
#define LOCALE_SABBREVDAYNAME1 0x00000031
#define LOCALE_SABBREVDAYNAME2 0x00000032
#define LOCALE_SABBREVDAYNAME3 0x00000033
#define LOCALE_SABBREVDAYNAME4 0x00000034
#define LOCALE_SABBREVDAYNAME5 0x00000035
#define LOCALE_SABBREVDAYNAME6 0x00000036
#define LOCALE_SABBREVDAYNAME7 0x00000037
#define LOCALE_SMONTHNAME1 0x00000038
#define LOCALE_SMONTHNAME2 0x00000039
#define LOCALE_SMONTHNAME3 0x0000003A
#define LOCALE_SMONTHNAME4 0x0000003B
#define LOCALE_SMONTHNAME5 0x0000003C
#define LOCALE_SMONTHNAME6 0x0000003D
#define LOCALE_SMONTHNAME7 0x0000003E
#define LOCALE_SMONTHNAME8 0x0000003F
#define LOCALE_SMONTHNAME9 0x00000040
#define LOCALE_SMONTHNAME10 0x00000041
#define LOCALE_SMONTHNAME11 0x00000042
#define LOCALE_SMONTHNAME12 0x00000043
#define LOCALE_SMONTHNAME13 0x0000100E
#define LOCALE_SABBREVMONTHNAME1 0x00000044
#define LOCALE_SABBREVMONTHNAME2 0x00000045
#define LOCALE_SABBREVMONTHNAME3 0x00000046
#define LOCALE_SABBREVMONTHNAME4 0x00000047
#define LOCALE_SABBREVMONTHNAME5 0x00000048
#define LOCALE_SABBREVMONTHNAME6 0x00000049
#define LOCALE_SABBREVMONTHNAME7 0x0000004A
#define LOCALE_SABBREVMONTHNAME8 0x0000004B
#define LOCALE_SABBREVMONTHNAME9 0x0000004C
#define LOCALE_SABBREVMONTHNAME10 0x0000004D
#define LOCALE_SABBREVMONTHNAME11 0x0000004E
#define LOCALE_SABBREVMONTHNAME12 0x0000004F
#define LOCALE_SABBREVMONTHNAME13 0x0000100F
#define LOCALE_SPOSITIVESIGN 0x00000050
#define LOCALE_SNEGATIVESIGN 0x00000051
#define LOCALE_IPOSSIGNPOSN 0x00000052
#define LOCALE_INEGSIGNPOSN 0x00000053
#define LOCALE_IPOSSYMPRECEDES 0x00000054
#define LOCALE_IPOSSEPBYSPACE 0x00000055
#define LOCALE_INEGSYMPRECEDES 0x00000056
#define LOCALE_INEGSEPBYSPACE 0x00000057
#define LOCALE_FONTSIGNATURE 0x00000058
#define TIME_NOMINUTESORSECONDS 0x00000001
#define TIME_NOSECONDS 0x00000002
#define TIME_NOTIMEMARKER 0x00000004
#define TIME_FORCE24HOURFORMAT 0x00000008
#define DATE_SHORTDATE 0x00000001
#define DATE_LONGDATE 0x00000002
#define DATE_USE_ALT_CALENDAR 0x00000004
#define CAL_ICALINTVALUE 0x00000001
#define CAL_SCALNAME 0x00000002
#define CAL_IYEAROFFSETRANGE 0x00000003
#define CAL_SERASTRING 0x00000004
#define CAL_SSHORTDATE 0x00000005
#define CAL_SLONGDATE 0x00000006
#define CAL_SDAYNAME1 0x00000007
#define CAL_SDAYNAME2 0x00000008
#define CAL_SDAYNAME3 0x00000009
#define CAL_SDAYNAME4 0x0000000a
#define CAL_SDAYNAME5 0x0000000b
#define CAL_SDAYNAME6 0x0000000c
#define CAL_SDAYNAME7 0x0000000d
#define CAL_SABBREVDAYNAME1 0x0000000e
#define CAL_SABBREVDAYNAME2 0x0000000f
#define CAL_SABBREVDAYNAME3 0x00000010
#define CAL_SABBREVDAYNAME4 0x00000011
#define CAL_SABBREVDAYNAME5 0x00000012
#define CAL_SABBREVDAYNAME6 0x00000013
#define CAL_SABBREVDAYNAME7 0x00000014
#define CAL_SMONTHNAME1 0x00000015
#define CAL_SMONTHNAME2 0x00000016
#define CAL_SMONTHNAME3 0x00000017
#define CAL_SMONTHNAME4 0x00000018
#define CAL_SMONTHNAME5 0x00000019
#define CAL_SMONTHNAME6 0x0000001a
#define CAL_SMONTHNAME7 0x0000001b
#define CAL_SMONTHNAME8 0x0000001c
#define CAL_SMONTHNAME9 0x0000001d
#define CAL_SMONTHNAME10 0x0000001e
#define CAL_SMONTHNAME11 0x0000001f
#define CAL_SMONTHNAME12 0x00000020
#define CAL_SMONTHNAME13 0x00000021
#define CAL_SABBREVMONTHNAME1 0x00000022
#define CAL_SABBREVMONTHNAME2 0x00000023
#define CAL_SABBREVMONTHNAME3 0x00000024
#define CAL_SABBREVMONTHNAME4 0x00000025
#define CAL_SABBREVMONTHNAME5 0x00000026
#define CAL_SABBREVMONTHNAME6 0x00000027
#define CAL_SABBREVMONTHNAME7 0x00000028
#define CAL_SABBREVMONTHNAME8 0x00000029
#define CAL_SABBREVMONTHNAME9 0x0000002a
#define CAL_SABBREVMONTHNAME10 0x0000002b
#define CAL_SABBREVMONTHNAME11 0x0000002c
#define CAL_SABBREVMONTHNAME12 0x0000002d
#define CAL_SABBREVMONTHNAME13 0x0000002e
#define ENUM_ALL_CALENDARS 0xffffffff
#define CAL_GREGORIAN 1
#define CAL_GREGORIAN_US 2
#define CAL_JAPAN 3
#define CAL_TAIWAN 4
#define CAL_KOREA 5
#define WC_NO_BEST_FIT_CHARS 0x00000400
#define MAP_EXPAND_LIGATURES 0x00002000
#define LCMAP_LINGUISTIC_CASING 0x01000000
#define LCMAP_SIMPLIFIED_CHINESE 0x02000000
#define LCMAP_TRADITIONAL_CHINESE 0x04000000
#define CSTR_LESS_THAN 1
#define CSTR_EQUAL 2
#define CSTR_GREATER_THAN 3
#define CP_THREAD_ACP 3
#define CP_SYMBOL 42
#define CP_UTF7 65000
#define CP_UTF8 65001
#define CTRY_ALBANIA 355
#define CTRY_ALGERIA 213
#define CTRY_ARGENTINA 54
#define CTRY_BELARUS 375
#define CTRY_BELIZE 501
#define CTRY_BOLIVIA 591
#define CTRY_BRUNEI_DARUSSALAM 673
#define CTRY_CARIBBEAN 1
#define CTRY_CHILE 56
#define CTRY_COLOMBIA 57
#define CTRY_COSTA_RICA 506
#define CTRY_DOMINICAN_REPUBLIC 1
#define CTRY_ECUADOR 593
#define CTRY_EGYPT 20
#define CTRY_EL_SALVADOR 503
#define CTRY_ESTONIA 372
#define CTRY_FAEROE_ISLANDS 298
#define CTRY_GUATEMALA 502
#define CTRY_HONDURAS 504
#define CTRY_INDIA 91
#define CTRY_INDONESIA 62
#define CTRY_IRAN 981
#define CTRY_IRAQ 964
#define CTRY_ISRAEL 972
#define CTRY_JAMAICA 1
#define CTRY_JORDAN 962
#define CTRY_KENYA 254
#define CTRY_KUWAIT 965
#define CTRY_LATVIA 371
#define CTRY_LEBANON 961
#define CTRY_LIBYA 218
#define CTRY_LIECHTENSTEIN 41
#define CTRY_LITHUANIA 370
#define CTRY_LUXEMBOURG 352
#define CTRY_MACAU 853
#define CTRY_MACEDONIA 389
#define CTRY_MALAYSIA 60
#define CTRY_MONACO 33
#define CTRY_MOROCCO 212
#define CTRY_NICARAGUA 505
#define CTRY_OMAN 968
#define CTRY_PAKISTAN 92
#define CTRY_PANAMA 507
#define CTRY_PARAGUAY 595
#define CTRY_PERU 51
#define CTRY_PHILIPPINES 63
#define CTRY_PUERTO_RICO 1
#define CTRY_QATAR 974
#define CTRY_SAUDI_ARABIA 966
#define CTRY_SERBIA 381
#define CTRY_SOUTH_AFRICA 27
#define CTRY_SYRIA 963
#define CTRY_THAILAND 66
#define CTRY_TRINIDAD_Y_TOBAGO 1
#define CTRY_TUNISIA 216
#define CTRY_UAE 971
#define CTRY_UKRAINE 380
#define CTRY_URUGUAY 598
#define CTRY_VENEZUELA 58
#define CTRY_VIET_NAM 84
#define CTRY_YEMEN 967
#define CTRY_ZIMBABWE 263
#define LOCALE_RETURN_NUMBER 0x20000000
#define LOCALE_IDEFAULTMACCODEPAGE 0x00001011
#define LOCALE_SISO639LANGNAME 0x00000059
#define LOCALE_SISO3166CTRYNAME 0x0000005A
#define LOCALE_IDEFAULTEBCDICCODEPAGE 0x00001012
#define LOCALE_IPAPERSIZE 0x0000100A
#define LOCALE_SENGCURRNAME 0x00001007
#define LOCALE_SNATIVECURRNAME 0x00001008
#define LOCALE_SYEARMONTH 0x00001006
#define LOCALE_SSORTNAME 0x00001013
#define LOCALE_IDIGITSUBSTITUTION 0x00001014
#define DATE_YEARMONTH 0x00000008
#define DATE_LTRREADING 0x00000010
#define DATE_RTLREADING 0x00000020
#define CAL_SYEARMONTH 0x0000002f
#define CAL_HIJRI 6
#define CAL_THAI 7
#define CAL_HEBREW 8
#define CAL_GREGORIAN_ME_FRENCH 9
#define CAL_GREGORIAN_ARABIC 10
#define CAL_GREGORIAN_XLIT_ENGLISH 11
#define CAL_GREGORIAN_XLIT_FRENCH 12
#define ANYSIZE_ARRAY 1
#define APPLICATION_ERROR_MASK 0x20000000
#define ERROR_SEVERITY_SUCCESS 0x00000000
#define ERROR_SEVERITY_INFORMATIONAL 0x40000000
#define ERROR_SEVERITY_WARNING 0x80000000
#define ERROR_SEVERITY_ERROR 0xC0000000
#define MINCHAR 0x80
#define MAXCHAR 0x7f
#define MINSHORT 0x8000
#define MAXSHORT 0x7fff
#define MINLONG 0x80000000
#define MAXBYTE 0xff
#define MAXWORD 0xffff
#define MAXDWORD 0xffffffff
#define LANG_NEUTRAL 0x00
#define LANG_INVARIANT 0x7f
#define LANG_AFRIKAANS 0x36
#define LANG_ALBANIAN 0x1c
#define LANG_ARABIC 0x01
#define LANG_ARMENIAN 0x2b
#define LANG_ASSAMESE 0x4d
#define LANG_AZERI 0x2c
#define LANG_BASQUE 0x2d
#define LANG_BELARUSIAN 0x23
#define LANG_BENGALI 0x45
#define LANG_BULGARIAN 0x02
#define LANG_CATALAN 0x03
#define LANG_CHINESE 0x04
#define LANG_CROATIAN 0x1a
#define LANG_CZECH 0x05
#define LANG_DANISH 0x06
#define LANG_DIVEHI 0x65
#define LANG_DUTCH 0x13
#define LANG_ENGLISH 0x09
#define LANG_ESTONIAN 0x25
#define LANG_FAEROESE 0x38
#define LANG_FARSI 0x29
#define LANG_FINNISH 0x0b
#define LANG_FRENCH 0x0c
#define LANG_GALICIAN 0x56
#define LANG_GEORGIAN 0x37
#define LANG_GERMAN 0x07
#define LANG_GREEK 0x08
#define LANG_GUJARATI 0x47
#define LANG_HEBREW 0x0d
#define LANG_HINDI 0x39
#define LANG_HUNGARIAN 0x0e
#define LANG_ICELANDIC 0x0f
#define LANG_INDONESIAN 0x21
#define LANG_ITALIAN 0x10
#define LANG_JAPANESE 0x11
#define LANG_KANNADA 0x4b
#define LANG_KASHMIRI 0x60
#define LANG_KAZAK 0x3f
#define LANG_KONKANI 0x57
#define LANG_KOREAN 0x12
#define LANG_KYRGYZ 0x40
#define LANG_LATVIAN 0x26
#define LANG_LITHUANIAN 0x27
#define LANG_MACEDONIAN 0x2f
#define LANG_MALAY 0x3e
#define LANG_MALAYALAM 0x4c
#define LANG_MANIPURI 0x58
#define LANG_MARATHI 0x4e
#define LANG_MONGOLIAN 0x50
#define LANG_NEPALI 0x61
#define LANG_NORWEGIAN 0x14
#define LANG_ORIYA 0x48
#define LANG_POLISH 0x15
#define LANG_PORTUGUESE 0x16
#define LANG_PUNJABI 0x46
#define LANG_ROMANIAN 0x18
#define LANG_RUSSIAN 0x19
#define LANG_SANSKRIT 0x4f
#define LANG_SERBIAN 0x1a
#define LANG_SINDHI 0x59
#define LANG_SLOVAK 0x1b
#define LANG_SLOVENIAN 0x24
#define LANG_SPANISH 0x0a
#define LANG_SWAHILI 0x41
#define LANG_SWEDISH 0x1d
#define LANG_SYRIAC 0x5a
#define LANG_TAMIL 0x49
#define LANG_TATAR 0x44
#define LANG_TELUGU 0x4a
#define LANG_THAI 0x1e
#define LANG_TURKISH 0x1f
#define LANG_UKRAINIAN 0x22
#define LANG_URDU 0x20
#define LANG_UZBEK 0x43
#define LANG_VIETNAMESE 0x2a
#define SUBLANG_NEUTRAL 0x00
#define SUBLANG_DEFAULT 0x01
#define SUBLANG_SYS_DEFAULT 0x02
#define SUBLANG_ARABIC_SAUDI_ARABIA 0x01
#define SUBLANG_ARABIC_IRAQ 0x02
#define SUBLANG_ARABIC_EGYPT 0x03
#define SUBLANG_ARABIC_LIBYA 0x04
#define SUBLANG_ARABIC_ALGERIA 0x05
#define SUBLANG_ARABIC_MOROCCO 0x06
#define SUBLANG_ARABIC_TUNISIA 0x07
#define SUBLANG_ARABIC_OMAN 0x08
#define SUBLANG_ARABIC_YEMEN 0x09
#define SUBLANG_ARABIC_SYRIA 0x0a
#define SUBLANG_ARABIC_JORDAN 0x0b
#define SUBLANG_ARABIC_LEBANON 0x0c
#define SUBLANG_ARABIC_KUWAIT 0x0d
#define SUBLANG_ARABIC_UAE 0x0e
#define SUBLANG_ARABIC_BAHRAIN 0x0f
#define SUBLANG_ARABIC_QATAR 0x10
#define SUBLANG_AZERI_LATIN 0x01
#define SUBLANG_AZERI_CYRILLIC 0x02
#define SUBLANG_CHINESE_TRADITIONAL 0x01
#define SUBLANG_CHINESE_SIMPLIFIED 0x02
#define SUBLANG_CHINESE_HONGKONG 0x03
#define SUBLANG_CHINESE_SINGAPORE 0x04
#define SUBLANG_CHINESE_MACAU 0x05
#define SUBLANG_DUTCH 0x01
#define SUBLANG_DUTCH_BELGIAN 0x02
#define SUBLANG_ENGLISH_US 0x01
#define SUBLANG_ENGLISH_UK 0x02
#define SUBLANG_ENGLISH_AUS 0x03
#define SUBLANG_ENGLISH_CAN 0x04
#define SUBLANG_ENGLISH_NZ 0x05
#define SUBLANG_ENGLISH_EIRE 0x06
#define SUBLANG_ENGLISH_SOUTH_AFRICA 0x07
#define SUBLANG_ENGLISH_JAMAICA 0x08
#define SUBLANG_ENGLISH_CARIBBEAN 0x09
#define SUBLANG_ENGLISH_BELIZE 0x0a
#define SUBLANG_ENGLISH_TRINIDAD 0x0b
#define SUBLANG_ENGLISH_ZIMBABWE 0x0c
#define SUBLANG_ENGLISH_PHILIPPINES 0x0d
#define SUBLANG_FRENCH 0x01
#define SUBLANG_FRENCH_BELGIAN 0x02
#define SUBLANG_FRENCH_CANADIAN 0x03
#define SUBLANG_FRENCH_SWISS 0x04
#define SUBLANG_FRENCH_LUXEMBOURG 0x05
#define SUBLANG_FRENCH_MONACO 0x06
#define SUBLANG_GERMAN 0x01
#define SUBLANG_GERMAN_SWISS 0x02
#define SUBLANG_GERMAN_AUSTRIAN 0x03
#define SUBLANG_GERMAN_LUXEMBOURG 0x04
#define SUBLANG_GERMAN_LIECHTENSTEIN 0x05
#define SUBLANG_ITALIAN 0x01
#define SUBLANG_ITALIAN_SWISS 0x02
#define SUBLANG_KASHMIRI_SASIA 0x02
#define SUBLANG_KASHMIRI_INDIA 0x02
#define SUBLANG_KOREAN 0x01
#define SUBLANG_LITHUANIAN 0x01
#define SUBLANG_MALAY_MALAYSIA 0x01
#define SUBLANG_MALAY_BRUNEI_DARUSSALAM 0x02
#define SUBLANG_NEPALI_INDIA 0x02
#define SUBLANG_NORWEGIAN_BOKMAL 0x01
#define SUBLANG_NORWEGIAN_NYNORSK 0x02
#define SUBLANG_PORTUGUESE 0x02
#define SUBLANG_PORTUGUESE_BRAZILIAN 0x01
#define SUBLANG_SERBIAN_LATIN 0x02
#define SUBLANG_SERBIAN_CYRILLIC 0x03
#define SUBLANG_SPANISH 0x01
#define SUBLANG_SPANISH_MEXICAN 0x02
#define SUBLANG_SPANISH_MODERN 0x03
#define SUBLANG_SPANISH_GUATEMALA 0x04
#define SUBLANG_SPANISH_COSTA_RICA 0x05
#define SUBLANG_SPANISH_PANAMA 0x06
#define SUBLANG_SPANISH_DOMINICAN_REPUBLIC 0x07
#define SUBLANG_SPANISH_VENEZUELA 0x08
#define SUBLANG_SPANISH_COLOMBIA 0x09
#define SUBLANG_SPANISH_PERU 0x0a
#define SUBLANG_SPANISH_ARGENTINA 0x0b
#define SUBLANG_SPANISH_ECUADOR 0x0c
#define SUBLANG_SPANISH_CHILE 0x0d
#define SUBLANG_SPANISH_URUGUAY 0x0e
#define SUBLANG_SPANISH_PARAGUAY 0x0f
#define SUBLANG_SPANISH_BOLIVIA 0x10
#define SUBLANG_SPANISH_EL_SALVADOR 0x11
#define SUBLANG_SPANISH_HONDURAS 0x12
#define SUBLANG_SPANISH_NICARAGUA 0x13
#define SUBLANG_SPANISH_PUERTO_RICO 0x14
#define SUBLANG_SWEDISH 0x01
#define SUBLANG_SWEDISH_FINLAND 0x02
#define SUBLANG_URDU_PAKISTAN 0x01
#define SUBLANG_URDU_INDIA 0x02
#define SUBLANG_UZBEK_LATIN 0x01
#define SUBLANG_UZBEK_CYRILLIC 0x02
#define SORT_DEFAULT 0x0
#define SORT_JAPANESE_XJIS 0x0
#define SORT_JAPANESE_UNICODE 0x1
#define SORT_CHINESE_BIG5 0x0
#define SORT_CHINESE_PRCP 0x0
#define SORT_CHINESE_UNICODE 0x1
#define SORT_CHINESE_PRC 0x2
#define SORT_CHINESE_BOPOMOFO 0x3
#define SORT_KOREAN_KSC 0x0
#define SORT_KOREAN_UNICODE 0x1
#define SORT_GERMAN_PHONE_BOOK 0x1
#define SORT_HUNGARIAN_DEFAULT 0x0
#define SORT_HUNGARIAN_TECHNICAL 0x1
#define SORT_GEORGIAN_TRADITIONAL 0x0
#define SORT_GEORGIAN_MODERN 0x1
#define NLS_VALID_LOCALE_MASK 0x000fffffU
#define LANG_SYSTEM_DEFAULT 0x0000002
#define LANG_USER_DEFAULT 0x0000001
#define LOCALE_SYSTEM_DEFAULT 0x800
#define LOCALE_USER_DEFAULT 0x400
#define LOCALE_NEUTRAL 0x0000
#define LOCALE_INVARIANT 0x007f
#define STATUS_NO_MEMORY DWORD (_CAST, 0xC0000017L)
#define MAXIMUM_WAIT_OBJECTS 64
#define MAXIMUM_SUSPEND_COUNT MAXCHAR
#define MAXIMUM_SUPPORTED_EXTENSION 512
#define SIZE_OF_80387_REGISTERS 80
#define CONTEXT_i386 0x00010000
#define CONTEXT_i486 0x00010000
#define CONTEXT_CONTROL 0x00010001L
#define CONTEXT_INTEGER 0x00010002L
#define CONTEXT_SEGMENTS 0x00010004L
#define CONTEXT_FLOATING_POINT 0x00010008L
#define CONTEXT_DEBUG_REGISTERS 0x00010010L
#define CONTEXT_FULL 0x00010007L
#define EXCEPTION_NONCONTINUABLE 0x1
#define EXCEPTION_MAXIMUM_PARAMETERS 15
#define PROCESS_TERMINATE 0x0001
#define PROCESS_CREATE_THREAD 0x0002
#define PROCESS_VM_OPERATION 0x0008
#define PROCESS_VM_READ 0x0010
#define PROCESS_VM_WRITE 0x0020
#define PROCESS_DUP_HANDLE 0x0040
#define PROCESS_CREATE_PROCESS 0x0080
#define PROCESS_SET_QUOTA 0x0100
#define PROCESS_SET_INFORMATION 0x0200
#define PROCESS_QUERY_INFORMATION 0x0400
#define PROCESS_ALL_ACCESS 0x001F0FFFl
#define THREAD_TERMINATE 0x0001
#define THREAD_SUSPEND_RESUME 0x0002
#define THREAD_GET_CONTEXT 0x0008
#define THREAD_SET_CONTEXT 0x0010
#define THREAD_SET_INFORMATION 0x0020
#define THREAD_QUERY_INFORMATION 0x0040
#define THREAD_SET_THREAD_TOKEN 0x0080
#define THREAD_IMPERSONATE 0x0100
#define THREAD_DIRECT_IMPERSONATION 0x0200
#define THREAD_ALL_ACCESS 0x001F03FFl
#define TLS_MINIMUM_AVAILABLE 64
#define EVENT_MODIFY_STATE 0x0002
#define EVENT_ALL_ACCESS 0x001F0003
#define SEMAPHORE_MODIFY_STATE 0x0002
#define SEMAPHORE_ALL_ACCESS 0x001F0003
#define TIME_ZONE_ID_UNKNOWN 0
#define TIME_ZONE_ID_STANDARD 1
#define TIME_ZONE_ID_DAYLIGHT 2
#define PROCESSOR_INTEL_386 386
#define PROCESSOR_INTEL_486 486
#define PROCESSOR_INTEL_PENTIUM 586
#define PROCESSOR_MIPS_R4000 4000
#define PROCESSOR_ALPHA_21064 21064
#define PROCESSOR_ARCHITECTURE_INTEL 0
#define PROCESSOR_ARCHITECTURE_MIPS 1
#define PROCESSOR_ARCHITECTURE_ALPHA 2
#define PROCESSOR_ARCHITECTURE_PPC 3
#define PROCESSOR_ARCHITECTURE_UNKNOWN 0xFFFF
#define SECTION_MAP_EXECUTE 0x0008
#define SECTION_EXTEND_SIZE 0x0010
#define PAGE_NOACCESS 0x01
#define PAGE_READONLY 0x02
#define PAGE_READWRITE 0x04
#define PAGE_WRITECOPY 0x08
#define PAGE_EXECUTE 0x10
#define PAGE_EXECUTE_READ 0x20
#define PAGE_EXECUTE_READWRITE 0x40
#define PAGE_EXECUTE_WRITECOPY 0x80
#define PAGE_GUARD 0x100
#define PAGE_NOCACHE 0x200
#define MEM_COMMIT 0x1000
#define MEM_RESERVE 0x2000
#define MEM_DECOMMIT 0x4000
#define MEM_RELEASE 0x8000
#define MEM_FREE 0x10000
#define MEM_PRIVATE 0x20000
#define MEM_MAPPED 0x40000
#define MEM_TOP_DOWN 0x100000
#define SEC_FILE 0x800000
#define SEC_IMAGE 0x1000000
#define SEC_RESERVE 0x4000000
#define SEC_COMMIT 0x8000000
#define SEC_NOCACHE 0x10000000
#define MEM_IMAGE SEC_IMAGE
#define FILE_READ_DATA 0x0001
#define FILE_LIST_DIRECTORY 0x0001
#define FILE_WRITE_DATA 0x0002
#define FILE_ADD_FILE 0x0002
#define FILE_APPEND_DATA 0x0004
#define FILE_ADD_SUBDIRECTORY 0x0004
#define FILE_CREATE_PIPE_INSTANCE 0x0004
#define FILE_READ_EA 0x0008
#define FILE_READ_PROPERTIES FILE_READ_EA
#define FILE_WRITE_EA 0x0010
#define FILE_WRITE_PROPERTIES FILE_WRITE_EA
#define FILE_EXECUTE 0x0020
#define FILE_TRAVERSE 0x0020
#define FILE_DELETE_CHILD 0x0040
#define FILE_READ_ATTRIBUTES 0x0080
#define FILE_WRITE_ATTRIBUTES 0x0100
#define FILE_ALL_ACCESS 0x001F01FFl
#define FILE_GENERIC_READ 0x00110089l
#define FILE_GENERIC_WRITE 0x00110116
#define FILE_GENERIC_EXECUTE 0x001f00A0
#define FILE_SHARE_READ 0x00000001
#define FILE_SHARE_WRITE 0x00000002
#define FILE_ATTRIBUTE_READONLY 0x00000001
#define FILE_ATTRIBUTE_HIDDEN 0x00000002
#define FILE_ATTRIBUTE_SYSTEM 0x00000004
#define FILE_ATTRIBUTE_DIRECTORY 0x00000010
#define FILE_ATTRIBUTE_ARCHIVE 0x00000020
#define FILE_ATTRIBUTE_NORMAL 0x00000080
#define FILE_ATTRIBUTE_TEMPORARY 0x00000100
#define FILE_ATTRIBUTE_COMPRESSED 0x00000800
#define FILE_NOTIFY_CHANGE_FILE_NAME 0x00000001
#define FILE_NOTIFY_CHANGE_DIR_NAME 0x00000002
#define FILE_NOTIFY_CHANGE_ATTRIBUTES 0x00000004
#define FILE_NOTIFY_CHANGE_SIZE 0x00000008
#define FILE_NOTIFY_CHANGE_LAST_WRITE 0x00000010
#define FILE_NOTIFY_CHANGE_SECURITY 0x00000100
#define MAILSLOT_NO_MESSAGE -1
#define MAILSLOT_WAIT_FOREVER -1
#define IO_COMPLETION_MODIFY_STATE 0x0002
#define IO_COMPLETION_ALL_ACCESS 0x001f0003l
#define DUPLICATE_CLOSE_SOURCE 0x00000001
#define DUPLICATE_SAME_ACCESS 0x00000002
//#define DELETE 0x00010000L
#define READ_CONTROL 0x00020000L
#define WRITE_DAC 0x00040000L
#define WRITE_OWNER 0x00080000L
#define SYNCHRONIZE 0x00100000L
#define STANDARD_RIGHTS_REQUIRED 0x000F0000L
#define STANDARD_RIGHTS_READ (READ_CONTROL)
#define STANDARD_RIGHTS_WRITE (READ_CONTROL)
#define STANDARD_RIGHTS_EXECUTE (READ_CONTROL)
#define STANDARD_RIGHTS_ALL 0x001F0000L
#define SPECIFIC_RIGHTS_ALL 0x0000FFFFL
#define ACCESS_SYSTEM_SECURITY 0x01000000L
#define MAXIMUM_ALLOWED 0x02000000L
#define GENERIC_READ 0x80000000L
#define GENERIC_WRITE 0x40000000L
#define GENERIC_EXECUTE 0x20000000L
#define GENERIC_ALL 0x10000000L
#define SID_REVISION 1
#define SID_MAX_SUB_AUTHORITIES 15
#define SID_RECOMMENDED_SUB_AUTHORITIES 1
#define SidTypeUser 1
#define SidTypeGroup 2
#define SidTypeDomain 3
#define SidTypeAlias 4
#define SidTypeWellKnownGroup 5
#define SidTypeDeletedAccount 6
#define SidTypeInvalid 7
#define SidTypeUnknown 8
#define SECURITY_NULL_RID 0x00000000L
#define SECURITY_WORLD_RID 0x00000000L
#define SECURITY_LOCAL_RID 0X00000000L
#define SECURITY_CREATOR_OWNER_RID 0x00000000L
#define SECURITY_CREATOR_GROUP_RID 0x00000001L
#define SECURITY_DIALUP_RID 0x00000001L
#define SECURITY_NETWORK_RID 0x00000002L
#define SECURITY_BATCH_RID 0x00000003L
#define SECURITY_INTERACTIVE_RID 0x00000004L
#define SECURITY_SERVICE_RID 0x00000006L
#define SECURITY_ANONYMOUS_LOGON_RID 0x00000007L
#define SECURITY_LOGON_IDS_RID 0x00000005L
#define SECURITY_LOGON_IDS_RID_COUNT 3L
#define SECURITY_LOCAL_SYSTEM_RID 0x00000012L
#define SECURITY_NT_NON_UNIQUE 0x00000015L
#define SECURITY_BUILTIN_DOMAIN_RID 0x00000020L
#define DOMAIN_USER_RID_ADMIN 0x000001F4L
#define DOMAIN_USER_RID_GUEST 0x000001F5L
#define DOMAIN_GROUP_RID_ADMINS 0x00000200L
#define DOMAIN_GROUP_RID_USERS 0x00000201L
#define DOMAIN_GROUP_RID_GUESTS 0x00000202L
#define DOMAIN_ALIAS_RID_ADMINS 0x00000220L
#define DOMAIN_ALIAS_RID_USERS 0x00000221L
#define DOMAIN_ALIAS_RID_GUESTS 0x00000222L
#define DOMAIN_ALIAS_RID_POWER_USERS 0x00000223L
#define DOMAIN_ALIAS_RID_ACCOUNT_OPS 0x00000224L
#define DOMAIN_ALIAS_RID_SYSTEM_OPS 0x00000225L
#define DOMAIN_ALIAS_RID_PRINT_OPS 0x00000226L
#define DOMAIN_ALIAS_RID_BACKUP_OPS 0x00000227L
#define DOMAIN_ALIAS_RID_REPLICATOR 0x00000228L
#define SE_GROUP_MANDATORY 0x00000001L
#define SE_GROUP_ENABLED_BY_DEFAULT 0x00000002L
#define SE_GROUP_ENABLED 0x00000004L
#define SE_GROUP_OWNER 0x00000008L
#define SE_GROUP_LOGON_ID 0xC0000000L
#define ACL_REVISION 2
#define ACL_REVISION1 1
#define ACL_REVISION2 2
#define ACCESS_ALLOWED_ACE_TYPE 0x0
#define ACCESS_DENIED_ACE_TYPE 0x1
#define SYSTEM_AUDIT_ACE_TYPE 0x2
#define SYSTEM_ALARM_ACE_TYPE 0x3
#define OBJECT_INHERIT_ACE 0x1
#define CONTAINER_INHERIT_ACE 0x2
#define NO_PROPAGATE_INHERIT_ACE 0x4
#define INHERIT_ONLY_ACE 0x8
#define VALID_INHERIT_FLAGS 0xF
#define SUCCESSFUL_ACCESS_ACE_FLAG 0x40
#define FAILED_ACCESS_ACE_FLAG 0x80
#define AclRevisionInformaton 1
#define AclSizeInformation 2
#define SECURITY_DESCRIPTOR_REVISION 1
#define SECURITY_DESCRIPTOR_REVISION1 1
#define SECURITY_DESCRIPTOR_MIN_LENGTH 20
#define SE_OWNER_DEFAULTED 0x0001
#define SE_GROUP_DEFAULTED 0x0002
#define SE_DACL_PRESENT 0x0004
#define SE_DACL_DEFAULTED 0x0008
#define SE_SACL_PRESENT 0x0010
#define SE_SACL_DEFAULTED 0x0020
#define SE_SELF_RELATIVE 0x8000
#define SE_PRIVILEGE_ENABLED_BY_DEFAULT 0x00000001
#define SE_PRIVILEGE_ENABLED 0x00000002
#define SE_PRIVILEGE_USED_FOR_ACCESS 0x80000000
#define PRIVILEGE_SET_ALL_NECESSARY 1
#define SE_CREATE_TOKEN_NAME "SeCreateTokenPrivilege"
#define SE_ASSIGNPRIMARYTOKEN_NAME "SeAssignPrimaryTokenPrivilege"
#define SE_LOCK_MEMORY_NAME "SeLockMemoryPrivilege"
#define SE_INCREASE_QUOTA_NAME "SeIncreaseQuotaPrivilege"
#define SE_UNSOLICITED_INPUT_NAME "SeUnsolicitedInputPrivilege"
#define SE_MACHINE_ACCOUNT_NAME "SeMachineAccountPrivilege"
#define SE_TCB_NAME "SeTcbPrivilege"
#define SE_SECURITY_NAME "SeSecurityPrivilege"
#define SE_TAKE_OWNERSHIP_NAME "SeTakeOwnershipPrivilege"
#define SE_LOAD_DRIVER_NAME "SeLoadDriverPrivilege"
#define SE_SYSTEM_PROFILE_NAME "SeSystemProfilePrivilege"
#define SE_SYSTEMTIME_NAME "SeSystemtimePrivilege"
#define SE_PROF_SINGLE_PROCESS_NAME "SeProfileSingleProcessPrivilege"
#define SE_INC_BASE_PRIORITY_NAME "SeIncreaseBasePriorityPrivilege"
#define SE_CREATE_PAGEFILE_NAME "SeCreatePagefilePrivilege"
#define SE_CREATE_PERMANENT_NAME "SeCreatePermanentPrivilege"
#define SE_BACKUP_NAME "SeBackupPrivilege"
#define SE_RESTORE_NAME "SeRestorePrivilege"
#define SE_SHUTDOWN_NAME "SeShutdownPrivilege"
#define SE_DEBUG_NAME "SeDebugPrivilege"
#define SE_AUDIT_NAME "SeAuditPrivilege"
#define SE_SYSTEM_ENVIRONMENT_NAME "SeSystemEnvironmentPrivilege"
#define SE_CHANGE_NOTIFY_NAME "SeChangeNotifyPrivilege"
#define SE_REMOTE_SHUTDOWN_NAME "SeRemoteShutdownPrivilege"
#define SecurityAnonymous 0
#define SecurityIdentification 1
#define SecurityImpersonation 2
#define SecurityDelegation 3
#define SECURITY_MAX_IMPERSONATION_LEVEL SecurityDelegation
#define DEFAULT_IMPERSONATION_LEVEL SecurityImpersonation
#define SECURITY_DYNAMIC_TRACKING TRUE
#define SECURITY_STATIC_TRACKING FALSE
#define TOKEN_ASSIGN_PRIMARY 0x0001
#define TOKEN_DUPLICATE 0x0002
#define TOKEN_IMPERSONATE 0x0004
#define TOKEN_QUERY 0x0008
#define TOKEN_QUERY_SOURCE 0x0010
#define TOKEN_ADJUST_PRIVILEGES 0x0020
#define TOKEN_ADJUST_GROUPS 0x0040
#define TOKEN_ADJUST_DEFAULT 0x0080
#define TOKEN_ALL_ACCESS 0X000F00FF
#define TOKEN_READ 0x00010008l
#define TOKEN_WRITE 0x000100E0l
#define TOKEN_EXECUTE (STANDARD_RIGHTS_EXECUTE)
#define TokenPrimary 1
#define TokenImpersonation 2
#define TokenUser 1
#define TokenGroups 2
#define TokenPrivileges 3
#define TokenOwner 4
#define TokenPrimaryGroup 5
#define TokenDefaultDacl 6
#define TokenSource 7
#define TokenType 8
#define TokenImpersonationLevel 9
#define TokenStatistics 10
#define TOKEN_SOURCE_LENGTH 8
#define OWNER_SECURITY_INFORMATION 0X00000001L
#define GROUP_SECURITY_INFORMATION 0X00000002L
#define DACL_SECURITY_INFORMATION 0X00000004L
#define SACL_SECURITY_INFORMATION 0X00000008L
#define IMAGE_DOS_SIGNATURE 0x5A4D
#define IMAGE_OS2_SIGNATURE 0x454E
#define IMAGE_OS2_SIGNATURE_LE 0x454C
#define IMAGE_VXD_SIGNATURE 0x454C
#define IMAGE_NT_SIGNATURE 0x00004550
#define IMAGE_SIZEOF_FILE_HEADER 20
#define IMAGE_FILE_RELOCS_STRIPPED 0x0001
#define IMAGE_FILE_EXECUTABLE_IMAGE 0x0002
#define IMAGE_FILE_LINE_NUMS_STRIPPED 0x0004
#define IMAGE_FILE_LOCAL_SYMS_STRIPPED 0x0008
#define IMAGE_FILE_AGGRESIVE_WS_TRIM 0x0010
#define IMAGE_FILE_LARGE_ADDRESS_AWARE 0x0020
#define IMAGE_FILE_BYTES_REVERSED_LO 0x0080
#define IMAGE_FILE_32BIT_MACHINE 0x0100
#define IMAGE_FILE_DEBUG_STRIPPED 0x0200
#define IMAGE_FILE_REMOVABLE_RUN_FROM_SWAP 0x0400
#define IMAGE_FILE_NET_RUN_FROM_SWAP 0x0800
#define IMAGE_FILE_SYSTEM 0x1000
#define IMAGE_FILE_DLL 0x2000
#define IMAGE_FILE_UP_SYSTEM_ONLY 0x4000
#define IMAGE_FILE_BYTES_REVERSED_HI 0x8000
#define IMAGE_FILE_MACHINE_UNKNOWN 0
#define IMAGE_FILE_MACHINE_I386 0x014c
#define IMAGE_FILE_MACHINE_R3000 0x0162
#define IMAGE_FILE_MACHINE_R4000 0x0166
#define IMAGE_FILE_MACHINE_R10000 0x0168
#define IMAGE_FILE_MACHINE_WCEMIPSV2 0x0169
#define IMAGE_FILE_MACHINE_ALPHA 0x0184
#define IMAGE_FILE_MACHINE_SH3 0x01a2
#define IMAGE_FILE_MACHINE_SH3DSP 0x01a3
#define IMAGE_FILE_MACHINE_SH3E 0x01a4
#define IMAGE_FILE_MACHINE_SH4 0x01a6
#define IMAGE_FILE_MACHINE_SH5 0x01a8
#define IMAGE_FILE_MACHINE_ARM 0x01c0
#define IMAGE_FILE_MACHINE_THUMB 0x01c2
#define IMAGE_FILE_MACHINE_AM33 0x01d3
#define IMAGE_FILE_MACHINE_POWERPC 0x01F0
#define IMAGE_FILE_MACHINE_POWERPCFP 0x01f1
#define IMAGE_FILE_MACHINE_IA64 0x0200
#define IMAGE_FILE_MACHINE_MIPS16 0x0266
#define IMAGE_FILE_MACHINE_ALPHA64 0x0284
#define IMAGE_FILE_MACHINE_MIPSFPU 0x0366
#define IMAGE_FILE_MACHINE_MIPSFPU16 0x0466
#define IMAGE_FILE_MACHINE_AXP64 IMAGE_FILE_MACHINE_ALPHA64
#define IMAGE_FILE_MACHINE_TRICORE 0x0520
#define IMAGE_FILE_MACHINE_CEF 0x0CEF
#define IMAGE_FILE_MACHINE_EBC 0x0EBC
#define IMAGE_FILE_MACHINE_AMD64 0x8664
#define IMAGE_FILE_MACHINE_M32R 0x9041
#define IMAGE_FILE_MACHINE_CEE 0xC0EE
#define IMAGE_NUMBEROF_DIRECTORY_ENTRIES 16
#define IMAGE_SIZEOF_ROM_OPTIONAL_HEADER 56
#define IMAGE_SIZEOF_STD_OPTIONAL_HEADER 28
#define IMAGE_SIZEOF_NT_OPTIONAL_HEADER 224
#define IMAGE_NT_OPTIONAL_HDR_MAGIC 0x10b
#define IMAGE_ROM_OPTIONAL_HDR_MAGIC 0x107
#define IMAGE_SUBSYSTEM_UNKNOWN 0
#define IMAGE_SUBSYSTEM_NATIVE 1
#define IMAGE_SUBSYSTEM_WINDOWS_GUI 2
#define IMAGE_SUBSYSTEM_WINDOWS_CUI 3
#define IMAGE_SUBSYSTEM_OS2_CUI 5
#define IMAGE_SUBSYSTEM_POSIX_CUI 7
#define IMAGE_DIRECTORY_ENTRY_EXPORT 0
#define IMAGE_DIRECTORY_ENTRY_IMPORT 1
#define IMAGE_DIRECTORY_ENTRY_RESOURCE 2
#define IMAGE_DIRECTORY_ENTRY_EXCEPTION 3
#define IMAGE_DIRECTORY_ENTRY_SECURITY 4
#define IMAGE_DIRECTORY_ENTRY_BASERELOC 5
#define IMAGE_DIRECTORY_ENTRY_DEBUG 6
#define IMAGE_DIRECTORY_ENTRY_COPYRIGHT 7
#define IMAGE_DIRECTORY_ENTRY_GLOBALPTR 8
#define IMAGE_DIRECTORY_ENTRY_TLS 9
#define IMAGE_DIRECTORY_ENTRY_LOAD_CONFIG 10
#define IMAGE_DIRECTORY_ENTRY_BOUND_IMPORT 11
#define IMAGE_DIRECTORY_ENTRY_IAT 12
#define IMAGE_SIZEOF_SHORT_NAME 8
#define IMAGE_SIZEOF_SECTION_HEADER 40
#define IMAGE_SCN_TYPE_NO_PAD 0x00000008
#define IMAGE_SCN_CNT_CODE 0x00000020
#define IMAGE_SCN_CNT_INITIALIZED_DATA 0x00000040
#define IMAGE_SCN_CNT_UNINITIALIZED_DATA 0x00000080
#define IMAGE_SCN_LNK_OTHER 0x00000100
#define IMAGE_SCN_LNK_INFO 0x00000200
#define IMAGE_SCN_LNK_REMOVE 0x00000800
#define IMAGE_SCN_LNK_COMDAT 0x00001000
#define IMAGE_SCN_MEM_FARDATA 0x00008000
#define IMAGE_SCN_MEM_PURGEABLE 0x00020000
#define IMAGE_SCN_MEM_16BIT 0x00020000
#define IMAGE_SCN_MEM_LOCKED 0x00040000
#define IMAGE_SCN_MEM_PRELOAD 0x00080000
#define IMAGE_SCN_ALIGN_1BYTES 0x00100000
#define IMAGE_SCN_ALIGN_2BYTES 0x00200000
#define IMAGE_SCN_ALIGN_4BYTES 0x00300000
#define IMAGE_SCN_ALIGN_8BYTES 0x00400000
#define IMAGE_SCN_ALIGN_16BYTES 0x00500000
#define IMAGE_SCN_ALIGN_32BYTES 0x00600000
#define IMAGE_SCN_ALIGN_64BYTES 0x00700000
#define IMAGE_SCN_LNK_NRELOC_OVFL 0x01000000
#define IMAGE_SCN_MEM_DISCARDABLE 0x02000000
#define IMAGE_SCN_MEM_NOT_CACHED 0x04000000
#define IMAGE_SCN_MEM_NOT_PAGED 0x08000000
#define IMAGE_SCN_MEM_SHARED 0x10000000
#define IMAGE_SCN_MEM_EXECUTE 0x20000000
#define IMAGE_SCN_MEM_READ 0x40000000
#define IMAGE_SCN_MEM_WRITE 0x80000000
#define IMAGE_SIZEOF_SYMBOL 18
#define IMAGE_SYM_ABSOLUTE -1
#define IMAGE_SYM_DEBUG -2
#define IMAGE_SYM_TYPE_NULL 0x0000
#define IMAGE_SYM_TYPE_VOID 0x0001
#define IMAGE_SYM_TYPE_CHAR 0x0002
#define IMAGE_SYM_TYPE_SHORT 0x0003
#define IMAGE_SYM_TYPE_INT 0x0004
#define IMAGE_SYM_TYPE_LONG 0x0005
#define IMAGE_SYM_TYPE_FLOAT 0x0006
#define IMAGE_SYM_TYPE_DOUBLE 0x0007
#define IMAGE_SYM_TYPE_STRUCT 0x0008
#define IMAGE_SYM_TYPE_UNION 0x0009
#define IMAGE_SYM_TYPE_ENUM 0x000A
#define IMAGE_SYM_TYPE_MOE 0x000B
#define IMAGE_SYM_TYPE_BYTE 0x000C
#define IMAGE_SYM_TYPE_WORD 0x000D
#define IMAGE_SYM_TYPE_UINT 0x000E
#define IMAGE_SYM_TYPE_DWORD 0x000F
#define IMAGE_SYM_TYPE_PCODE 0x8000
#define IMAGE_SYM_DTYPE_NULL 0
#define IMAGE_SYM_DTYPE_POINTER 1
#define IMAGE_SYM_DTYPE_FUNCTION 2
#define IMAGE_SYM_DTYPE_ARRAY 3
#define IMAGE_SYM_CLASS_END_OF_FUNCTION -1
#define IMAGE_SYM_CLASS_NULL 0x0000
#define IMAGE_SYM_CLASS_AUTOMATIC 0x0001
#define IMAGE_SYM_CLASS_EXTERNAL 0x0002
#define IMAGE_SYM_CLASS_STATIC 0x0003
#define IMAGE_SYM_CLASS_REGISTER 0x0004
#define IMAGE_SYM_CLASS_EXTERNAL_DEF 0x0005
#define IMAGE_SYM_CLASS_LABEL 0x0006
#define IMAGE_SYM_CLASS_UNDEFINED_LABEL 0x0007
#define IMAGE_SYM_CLASS_MEMBER_OF_STRUCT 0x0008
#define IMAGE_SYM_CLASS_ARGUMENT 0x0009
#define IMAGE_SYM_CLASS_STRUCT_TAG 0x000A
#define IMAGE_SYM_CLASS_MEMBER_OF_UNION 0x000B
#define IMAGE_SYM_CLASS_UNION_TAG 0x000C
#define IMAGE_SYM_CLASS_TYPE_DEFINITION 0x000D
#define IMAGE_SYM_CLASS_UNDEFINED_STATIC 0x000E
#define IMAGE_SYM_CLASS_ENUM_TAG 0x000F
#define IMAGE_SYM_CLASS_MEMBER_OF_ENUM 0x0010
#define IMAGE_SYM_CLASS_REGISTER_PARAM 0x0011
#define IMAGE_SYM_CLASS_BIT_FIELD 0x0012
#define IMAGE_SYM_CLASS_FAR_EXTERNAL 0x0044
#define IMAGE_SYM_CLASS_BLOCK 0x0064
#define IMAGE_SYM_CLASS_FUNCTION 0x0065
#define IMAGE_SYM_CLASS_END_OF_STRUCT 0x0066
#define IMAGE_SYM_CLASS_FILE 0x0067
#define IMAGE_SYM_CLASS_SECTION 0x0068
#define IMAGE_SYM_CLASS_WEAK_EXTERNAL 0x0069
#define N_BTMASK 0x000F
#define N_TMASK 0x0030
#define N_TMASK1 0x00C0
#define N_TMASK2 0x00F0
#define N_BTSHFT 4
#define N_TSHIFT 2
#define IMAGE_SIZEOF_AUX_SYMBOL 18
#define IMAGE_COMDAT_SELECT_NODUPLICATES 1
#define IMAGE_COMDAT_SELECT_ANY 2
#define IMAGE_COMDAT_SELECT_SAME_SIZE 3
#define IMAGE_COMDAT_SELECT_EXACT_MATCH 4
#define IMAGE_COMDAT_SELECT_ASSOCIATIVE 5
#define IMAGE_COMDAT_SELECT_LARGEST 6
#define IMAGE_COMDAT_SELECT_NEWEST 7
#define IMAGE_WEAK_EXTERN_SEARCH_NOLIBRARY 1
#define IMAGE_WEAK_EXTERN_SEARCH_LIBRARY 2
#define IMAGE_WEAK_EXTERN_SEARCH_ALIAS 3
#define IMAGE_SIZEOF_RELOCATION 10
#define IMAGE_REL_I386_ABSOLUTE 0x0000
#define IMAGE_REL_I386_DIR16 0x0001
#define IMAGE_REL_I386_REL16 0x0002
#define IMAGE_REL_I386_DIR32 0x0006
#define IMAGE_REL_I386_DIR32NB 0x0007
#define IMAGE_REL_I386_SEG12 0x0009
#define IMAGE_REL_I386_SECTION 0x000A
#define IMAGE_REL_I386_SECREL 0x000B
#define IMAGE_REL_I386_REL32 0x0014
#define IMAGE_REL_MIPS_ABSOLUTE 0x0000
#define IMAGE_REL_MIPS_REFHALF 0x0001
#define IMAGE_REL_MIPS_REFWORD 0x0002
#define IMAGE_REL_MIPS_JMPADDR 0x0003
#define IMAGE_REL_MIPS_REFHI 0x0004
#define IMAGE_REL_MIPS_REFLO 0x0005
#define IMAGE_REL_MIPS_GPREL 0x0006
#define IMAGE_REL_MIPS_LITERAL 0x0007
#define IMAGE_REL_MIPS_SECTION 0x000A
#define IMAGE_REL_MIPS_SECREL 0x000B
#define IMAGE_REL_MIPS_SECRELLO 0x000C
#define IMAGE_REL_MIPS_SECRELHI 0x000D
#define IMAGE_REL_MIPS_REFWORDNB 0x0022
#define IMAGE_REL_MIPS_PAIR 0x0025
#define IMAGE_REL_ALPHA_ABSOLUTE 0x0000
#define IMAGE_REL_ALPHA_REFLONG 0x0001
#define IMAGE_REL_ALPHA_REFQUAD 0x0002
#define IMAGE_REL_ALPHA_GPREL32 0x0003
#define IMAGE_REL_ALPHA_LITERAL 0x0004
#define IMAGE_REL_ALPHA_LITUSE 0x0005
#define IMAGE_REL_ALPHA_GPDISP 0x0006
#define IMAGE_REL_ALPHA_BRADDR 0x0007
#define IMAGE_REL_ALPHA_HINT 0x0008
#define IMAGE_REL_ALPHA_INLINE_REFLONG 0x0009
#define IMAGE_REL_ALPHA_REFHI 0x000A
#define IMAGE_REL_ALPHA_REFLO 0x000B
#define IMAGE_REL_ALPHA_PAIR 0x000C
#define IMAGE_REL_ALPHA_MATCH 0x000D
#define IMAGE_REL_ALPHA_SECTION 0x000E
#define IMAGE_REL_ALPHA_SECREL 0x000F
#define IMAGE_REL_ALPHA_REFLONGNB 0x0010
#define IMAGE_REL_ALPHA_SECRELLO 0x0011
#define IMAGE_REL_ALPHA_SECRELHI 0x0012
#define IMAGE_REL_PPC_ABSOLUTE 0x0000
#define IMAGE_REL_PPC_ADDR64 0x0001
#define IMAGE_REL_PPC_ADDR32 0x0002
#define IMAGE_REL_PPC_ADDR24 0x0003
#define IMAGE_REL_PPC_ADDR16 0x0004
#define IMAGE_REL_PPC_ADDR14 0x0005
#define IMAGE_REL_PPC_REL24 0x0006
#define IMAGE_REL_PPC_REL14 0x0007
#define IMAGE_REL_PPC_TOCREL16 0x0008
#define IMAGE_REL_PPC_TOCREL14 0x0009
#define IMAGE_REL_PPC_ADDR32NB 0x000A
#define IMAGE_REL_PPC_SECREL 0x000B
#define IMAGE_REL_PPC_SECTION 0x000C
#define IMAGE_REL_PPC_IFGLUE 0x000D
#define IMAGE_REL_PPC_IMGLUE 0x000E
#define IMAGE_REL_PPC_SECREL16 0x000F
#define IMAGE_REL_PPC_REFHI 0x0010
#define IMAGE_REL_PPC_REFLO 0x0011
#define IMAGE_REL_PPC_PAIR 0x0012
#define IMAGE_REL_PPC_TYPEMASK 0x00FF
#define IMAGE_REL_PPC_NEG 0x0100
#define IMAGE_REL_PPC_BRTAKEN 0x0200
#define IMAGE_REL_PPC_BRNTAKEN 0x0400
#define IMAGE_REL_PPC_TOCDEFN 0x0800
#define IMAGE_SIZEOF_BASE_RELOCATION 8
#define IMAGE_REL_BASED_ABSOLUTE 0
#define IMAGE_REL_BASED_HIGH 1
#define IMAGE_REL_BASED_LOW 2
#define IMAGE_REL_BASED_HIGHLOW 3
#define IMAGE_REL_BASED_HIGHADJ 4
#define IMAGE_REL_BASED_MIPS_JMPADDR 5
#define IMAGE_SIZEOF_LINENUMBER 6
#define IMAGE_ARCHIVE_START_SIZE 8
#define IMAGE_SIZEOF_ARCHIVE_MEMBER_HDR 60
#define IMAGE_ORDINAL_FLAG 0x80000000
#define IMAGE_RESOURCE_NAME_IS_STRING 0x80000000
#define IMAGE_RESOURCE_DATA_IS_DIRECTORY 0x80000000
#define IMAGE_DEBUG_TYPE_UNKNOWN 0
#define IMAGE_DEBUG_TYPE_COFF 1
#define IMAGE_DEBUG_TYPE_CODEVIEW 2
#define IMAGE_DEBUG_TYPE_FPO 3
#define IMAGE_DEBUG_TYPE_MISC 4
#define IMAGE_DEBUG_TYPE_EXCEPTION 5
#define IMAGE_DEBUG_TYPE_FIXUP 6
#define IMAGE_DEBUG_TYPE_OMAP_TO_SRC 7
#define IMAGE_DEBUG_TYPE_OMAP_FROM_SRC 8
#define FRAME_FPO 0
#define FRAME_TRAP 1
#define FRAME_TSS 2
#define FRAME_NONFPO 3
#define SIZEOF_RFPO_DATA 16
#define IMAGE_DEBUG_MISC_EXENAME 1
#define IMAGE_SEPARATE_DEBUG_SIGNATURE 0x4944
#define NON_PAGED_DEBUG_SIGNATURE 0x494E
#define IMAGE_SEPARATE_DEBUG_FLAGS_MASK 0x8000
#define IMAGE_SEPARATE_DEBUG_MISMATCH 0x8000
#define HEAP_NO_SERIALIZE 0x00000001
#define HEAP_GROWABLE 0x00000002
#define HEAP_GENERATE_EXCEPTIONS 0x00000004
#define HEAP_ZERO_MEMORY 0x00000008
#define HEAP_REALLOC_IN_PLACE_ONLY 0x00000010
#define HEAP_TAIL_CHECKING_ENABLED 0x00000020
#define HEAP_FREE_CHECKING_ENABLED 0x00000040
#define HEAP_DISABLE_COALESCE_ON_FREE 0x00000080
#define HEAP_CREATE_ALIGN_16 0x00010000
#define HEAP_CREATE_ENABLE_TRACING 0x00020000
#define HEAP_MAXIMUM_TAG 0x0FFF
#define HEAP_PSEUDO_TAG_FLAG 0x8000
#define HEAP_TAG_SHIFT 16
#define IS_TEXT_UNICODE_ASCII16 0x0001
#define IS_TEXT_UNICODE_REVERSE_ASCII16 0x0010
#define IS_TEXT_UNICODE_STATISTICS 0x0002
#define IS_TEXT_UNICODE_REVERSE_STATISTICS 0x0020
#define IS_TEXT_UNICODE_CONTROLS 0x0004
#define IS_TEXT_UNICODE_REVERSE_CONTROLS 0x0040
#define IS_TEXT_UNICODE_SIGNATURE 0x0008
#define IS_TEXT_UNICODE_REVERSE_SIGNATURE 0x0080
#define IS_TEXT_UNICODE_ILLEGAL_CHARS 0x0100
#define IS_TEXT_UNICODE_ODD_LENGTH 0x0200
#define IS_TEXT_UNICODE_DBCS_LEADBYTE 0x0400
#define IS_TEXT_UNICODE_NULL_BYTES 0x1000
#define IS_TEXT_UNICODE_UNICODE_MASK 0x000F
#define IS_TEXT_UNICODE_REVERSE_MASK 0x00F0
#define IS_TEXT_UNICODE_NOT_UNICODE_MASK 0x0F00
#define IS_TEXT_UNICODE_NOT_ASCII_MASK 0xF000
#define COMPRESSION_FORMAT_NONE (0x0000)
#define COMPRESSION_FORMAT_DEFAULT (0x0001)
#define COMPRESSION_FORMAT_LZNT1 (0x0002)
#define COMPRESSION_ENGINE_STANDARD (0x0000)
#define COMPRESSION_ENGINE_MAXIMUM (0x0100)
#define MESSAGE_RESOURCE_UNICODE 0x0001
#define RTL_CRITSECT_TYPE 0
#define RTL_RESOURCE_TYPE 1
#define DLL_PROCESS_ATTACH 1
#define DLL_THREAD_ATTACH 2
#define DLL_THREAD_DETACH 3
#define DLL_PROCESS_DETACH 0
#define EVENTLOG_SEQUENTIAL_READ 0X0001
#define EVENTLOG_SEEK_READ 0X0002
#define EVENTLOG_FORWARDS_READ 0X0004
#define EVENTLOG_BACKWARDS_READ 0X0008
#define EVENTLOG_SUCCESS 0X0000
#define EVENTLOG_ERROR_TYPE 0x0001
#define EVENTLOG_WARNING_TYPE 0x0002
#define EVENTLOG_INFORMATION_TYPE 0x0004
#define EVENTLOG_AUDIT_SUCCESS 0x0008
#define EVENTLOG_AUDIT_FAILURE 0x0010
#define EVENTLOG_START_PAIRED_EVENT 0x0001
#define EVENTLOG_END_PAIRED_EVENT 0x0002
#define EVENTLOG_END_ALL_PAIRED_EVENTS 0x0004
#define EVENTLOG_PAIRED_EVENT_ACTIVE 0x0008
#define EVENTLOG_PAIRED_EVENT_INACTIVE 0x0010
#define DBG_CONTINUE DWORD(_CAST,0x00010002)
#define DBG_TERMINATE_THREAD DWORD(_CAST,0x40010003)
#define DBG_TERMINATE_PROCESS DWORD(_CAST,0x40010004)
#define DBG_CONTROL_C DWORD(_CAST,0x40010005)
#define DBG_CONTROL_BREAK DWORD(_CAST,0x40010008)
#define DBG_EXCEPTION_NOT_HANDLED DWORD(_CAST,0x80010001)
#define KEY_QUERY_VALUE 0x0001
#define KEY_SET_VALUE 0x0002
#define KEY_CREATE_SUB_KEY 0x0004
#define KEY_ENUMERATE_SUB_KEYS 0x0008
#define KEY_NOTIFY 0x0010
#define KEY_CREATE_LINK 0x0020
#define KEY_WRITE 0x00020006U
#define KEY_READ 0x00020019U
#define KEY_ALL_ACCESS 0x000F003FU
#define REG_OPTION_RESERVED 0x00000000L
#define REG_OPTION_NON_VOLATILE 0x00000000L
#define REG_OPTION_VOLATILE 0x00000001L
#define REG_OPTION_CREATE_LINK 0x00000002L
#define REG_OPTION_BACKUP_RESTORE 0x00000004L
#define REG_LEGAL_OPTION 0x00000007L
#define REG_CREATED_NEW_KEY 0x00000001L
#define REG_OPENED_EXISTING_KEY 0x00000002L
#define REG_WHOLE_HIVE_VOLATILE 0x00000001L
#define REG_REFRESH_HIVE 0x00000002L
#define REG_NOTIFY_CHANGE_NAME 0x00000001L
#define REG_NOTIFY_CHANGE_ATTRIBUTES 0x00000002L
#define REG_NOTIFY_CHANGE_LAST_SET 0x00000004L
#define REG_NOTIFY_CHANGE_SECURITY 0x00000008L
#define REG_LEGAL_CHANGE_FILTER 0x0000000Fl
#define REG_NONE 0
#define REG_SZ 1
#define REG_EXPAND_SZ 2
#define REG_BINARY 3
#define REG_DWORD 4
#define REG_DWORD_LITTLE_ENDIAN 4
#define REG_DWORD_BIG_ENDIAN 5
#define REG_LINK 6
#define REG_MULTI_SZ 7
#define REG_RESOURCE_LIST 8
#define REG_FULL_RESOURCE_DESCRIPTOR 9
#define REG_RESOURCE_REQUIREMENTS_LIST 10
#define SERVICE_KERNEL_DRIVER 0x00000001
#define SERVICE_FILE_SYSTEM_DRIVER 0x00000002
#define SERVICE_ADAPTER 0x00000004
#define SERVICE_RECOGNIZER_DRIVER 0x00000008
#define SERVICE_DRIVER 0x0000000B
#define SERVICE_WIN32_OWN_PROCESS 0x00000010
#define SERVICE_WIN32_SHARE_PROCESS 0x00000020
#define SERVICE_WIN32 0x00000030L
#define SERVICE_INTERACTIVE_PROCESS 0x00000100
#define SERVICE_TYPE_ALL 0x0000013Fl
#define SERVICE_BOOT_START 0x00000000
#define SERVICE_SYSTEM_START 0x00000001
#define SERVICE_AUTO_START 0x00000002
#define SERVICE_DEMAND_START 0x00000003
#define SERVICE_DISABLED 0x00000004
#define SERVICE_ERROR_IGNORE 0x00000000
#define SERVICE_ERROR_NORMAL 0x00000001
#define SERVICE_ERROR_SEVERE 0x00000002
#define SERVICE_ERROR_CRITICAL 0x00000003
#define DriverType 0x00000001
#define FileSystemType 0x00000002
#define Win32ServiceOwnProcess 0x00000010
#define win32ServiceShareProcess 0x00000020
#define AdapterTyper 0x00000004
#define Recongnizertype 0x00000008
#define BootLoad 0x00000000
#define SystemLoad 0x00000001
#define AutoLoad 0x00000002
#define DemandLoad 0x00000003
#define DisableLoad 0x00000004
#define IgnoreError 0x00000000
#define NormalError 0x00000001
#define SevereError 0x00000002
#define CriticalError 0x00000003
#define TAPE_ERASE_SHORT 0L
#define TAPE_ERASE_LONG 1L
#define TAPE_LOAD 0L
#define TAPE_UNLOAD 1L
#define TAPE_TENSION 2L
#define TAPE_LOCK 3L
#define TAPE_UNLOCK 4L
#define TAPE_FORMAT 5L
#define TAPE_SETMARKS 0L
#define TAPE_FILEMARKS 1L
#define TAPE_SHORT_FILEMARKS 2L
#define TAPE_LONG_FILEMARKS 3L
#define TAPE_ABSOLUTE_POSITION 0L
#define TAPE_LOGICAL_POSITION 1L
#define TAPE_PSEUDO_LOGICAL_POSITION 2L
#define TAPE_REWIND 0L
#define TAPE_ABSOLUTE_BLOCK 1L
#define TAPE_LOGICAL_BLOCK 2L
#define TAPE_PSEUDO_LOGICAL_BLOCK 3L
#define TAPE_SPACE_END_OF_DATA 4L
#define TAPE_SPACE_RELATIVE_BLOCKS 5L
#define TAPE_SPACE_FILEMARKS 6L
#define TAPE_SPACE_SEQUENTIAL_FMKS 7L
#define TAPE_SPACE_SETMARKS 8L
#define TAPE_SPACE_SEQUENTIAL_SMKS 9L
#define TAPE_DRIVE_FIXED 0x00000001
#define TAPE_DRIVE_SELECT 0x00000002
#define TAPE_DRIVE_INITIATOR 0x00000004
#define TAPE_DRIVE_ERASE_SHORT 0x00000010
#define TAPE_DRIVE_ERASE_LONG 0x00000020
#define TAPE_DRIVE_ERASE_BOP_ONLY 0x00000040
#define TAPE_DRIVE_ERASE_IMMEDIATE 0x00000080
#define TAPE_DRIVE_TAPE_CAPACITY 0x00000100
#define TAPE_DRIVE_TAPE_REMAINING 0x00000200
#define TAPE_DRIVE_FIXED_BLOCK 0x00000400
#define TAPE_DRIVE_VARIABLE_BLOCK 0x00000800
#define TAPE_DRIVE_WRITE_PROTECT 0x00001000
#define TAPE_DRIVE_EOT_WZ_SIZE 0x00002000
#define TAPE_DRIVE_ECC 0x00010000
#define TAPE_DRIVE_COMPRESSION 0x00020000
#define TAPE_DRIVE_PADDING 0x00040000
#define TAPE_DRIVE_REPORT_SMKS 0x00080000
#define TAPE_DRIVE_GET_ABSOLUTE_BLK 0x00100000
#define TAPE_DRIVE_GET_LOGICAL_BLK 0x00200000
#define TAPE_DRIVE_SET_EOT_WZ_SIZE 0x00400000
#define TAPE_DRIVE_RESERVED_BIT 0x80000000
#define TAPE_DRIVE_LOAD_UNLOAD 0x80000001
#define TAPE_DRIVE_TENSION 0x80000002
#define TAPE_DRIVE_LOCK_UNLOCK 0x80000004
#define TAPE_DRIVE_REWIND_IMMEDIATE 0x80000008
#define TAPE_DRIVE_SET_BLOCK_SIZE 0x80000010
#define TAPE_DRIVE_LOAD_UNLD_IMMED 0x80000020
#define TAPE_DRIVE_TENSION_IMMED 0x80000040
#define TAPE_DRIVE_LOCK_UNLK_IMMED 0x80000080
#define TAPE_DRIVE_SET_ECC 0x80000100
#define TAPE_DRIVE_SET_COMPRESSION 0x80000200
#define TAPE_DRIVE_SET_PADDING 0x80000400
#define TAPE_DRIVE_SET_REPORT_SMKS 0x80000800
#define TAPE_DRIVE_ABSOLUTE_BLK 0x80001000
#define TAPE_DRIVE_ABS_BLK_IMMED 0x80002000
#define TAPE_DRIVE_LOGICAL_BLK 0x80004000
#define TAPE_DRIVE_LOG_BLK_IMMED 0x80008000
#define TAPE_DRIVE_END_OF_DATA 0x80010000
#define TAPE_DRIVE_RELATIVE_BLKS 0x80020000
#define TAPE_DRIVE_FILEMARKS 0x80040000
#define TAPE_DRIVE_SEQUENTIAL_FMKS 0x80080000
#define TAPE_DRIVE_SETMARKS 0x80100000
#define TAPE_DRIVE_SEQUENTIAL_SMKS 0x80200000
#define TAPE_DRIVE_REVERSE_POSITION 0x80400000
#define TAPE_DRIVE_SPACE_IMMEDIATE 0x80800000
#define TAPE_DRIVE_WRITE_SETMARKS 0x81000000
#define TAPE_DRIVE_WRITE_FILEMARKS 0x82000000
#define TAPE_DRIVE_WRITE_SHORT_FMKS 0x84000000
#define TAPE_DRIVE_WRITE_LONG_FMKS 0x88000000
#define TAPE_DRIVE_WRITE_MARK_IMMED 0x90000000
#define TAPE_DRIVE_FORMAT 0xA0000000
#define TAPE_DRIVE_FORMAT_IMMEDIATE 0xC0000000
#define TAPE_DRIVE_HIGH_FEATURES 0x80000000
#define TAPE_FIXED_PARTITIONS 0L
#define TAPE_SELECT_PARTITIONS 1L
#define TAPE_INITIATOR_PARTITIONS 2L
#define WT_EXECUTEDEFAULT 0x00000000
#define WT_EXECUTEINIOTHREAD 0x00000001
#define WT_EXECUTEINUITHREAD 0x00000002
#define WT_EXECUTEINWAITTHREAD 0x00000004
#define WT_EXECUTEDELETEWAIT 0x00000008
#define WT_EXECUTEINLONGTHREAD 0x00000010
#define IMAGE_SYM_UNDEFINED SHORTINT(_CAST,0)
#define PERF_DATA_VERSION 1
#define PERF_DATA_REVISION 1
#define PERF_NO_INSTANCES -1
#define PERF_SIZE_DWORD 0x00000000
#define PERF_SIZE_LARGE 0x00000100
#define PERF_SIZE_ZERO 0x00000200
#define PERF_SIZE_VARIABLE_LEN 0x00000300
#define PERF_TYPE_NUMBER 0x00000000
#define PERF_TYPE_COUNTER 0x00000400
#define PERF_TYPE_TEXT 0x00000800
#define PERF_TYPE_ZERO 0x00000C00
#define PERF_NUMBER_HEX 0x00000000
#define PERF_NUMBER_DECIMAL 0x00010000
#define PERF_NUMBER_DEC_1000 0x00020000
#define PERF_COUNTER_VALUE 0x00000000
#define PERF_COUNTER_RATE 0x00010000
#define PERF_COUNTER_FRACTION 0x00020000
#define PERF_COUNTER_BASE 0x00030000
#define PERF_COUNTER_ELAPSED 0x00040000
#define PERF_COUNTER_QUEUELEN 0x00050000
#define PERF_COUNTER_HISTOGRAM 0x00060000
#define PERF_COUNTER_PRECISION 0x00070000
#define PERF_TEXT_UNICODE 0x00000000
#define PERF_TEXT_ASCII 0x00010000
#define PERF_TIMER_TICK 0x00000000
#define PERF_TIMER_100NS 0x00100000
#define PERF_OBJECT_TIMER 0x00200000
#define PERF_DELTA_COUNTER 0x00400000
#define PERF_DELTA_BASE 0x00800000
#define PERF_INVERSE_COUNTER 0x01000000
#define PERF_MULTI_COUNTER 0x02000000
#define PERF_DISPLAY_NO_SUFFIX 0x00000000
#define PERF_DISPLAY_PER_SEC 0x10000000
#define PERF_DISPLAY_PERCENT 0x20000000
#define PERF_DISPLAY_SECONDS 0x30000000
#define PERF_DISPLAY_NOSHOW 0x40000000
#define PERF_COUNTER_COUNTER 0x10410400
#define PERF_COUNTER_TIMER 0x10410500
#define PERF_COUNTER_QUEUELEN_TYPE 0x00450400
#define PERF_COUNTER_BULK_COUNT 0x10410500
#define PERF_COUNTER_TEXT 0x00000B00
#define PERF_COUNTER_RAWCOUNT 0x00010000
#define PERF_COUNTER_LARGE_RAWCOUNT 0x00010100
#define PERF_COUNTER_RAWCOUNT_HEX 0x00000000
#define PERF_COUNTER_LARGE_RAWCOUNT_HEX 0x00000100
#define PERF_SAMPLE_FRACTION 0x20c20400
#define PERF_SAMPLE_COUNTER 0x00410400
#define PERF_COUNTER_NODATA 0x40000200
#define PERF_COUNTER_TIMER_INV 0x21410500
#define PERF_SAMPLE_BASE 0x40030401
#define PERF_AVERAGE_TIMER 0x30020400
#define PERF_AVERAGE_BASE 0x40030402
#define PERF_AVERAGE_BULK 0x4020500
#define PERF_100NSEC_TIMER 0x20510500
#define PERF_100NSEC_TIMER_INV 0x21500500
#define PERF_COUNTER_MULTI_TIMER 0x22410500
#define PERF_COUNTER_MULTI_TIMER_INV 0x23410500
#define PERF_COUNTER_MULTI_BASE 0x42030500
#define PERF_100NSEC_MULTI_TIMER 0x22510500
#define PERF_100NSEC_MULTI_TIMER_INV 0x23510500
#define PERF_RAW_FRACTION 0x20020400
#define PERF_RAW_BASE 0x40030403
#define PERF_ELAPSED_TIME 0x30240500
#define PERF_COUNTER_HISTOGRAM_TYPE 0x80000000
#define PERF_DETAIL_NOVICE 100
#define PERF_DETAIL_ADVANCED 200
#define PERF_DETAIL_EXPERT 300
#define PERF_DETAIL_WIZARD 400
#define PERF_NO_UNIQUE_ID -1
#define PERF_QUERY_OBJECTS 0x80000000L
#define PERF_QUERY_GLOBAL 0x80000001L
#define PERF_QUERY_COSTLY 0x80000002L
#define WINPERF_LOG_NONE 0
#define WINPERF_LOG_USER 1
#define WINPERF_LOG_DEBUG 2
#define WINPERF_LOG_VERBOSE 3
#define RRF_RT_REG_NONE 0x00000001
#define RRF_RT_REG_SZ 0x00000002
#define RRF_RT_REG_EXPAND_SZ 0x00000004
#define RRF_RT_REG_BINARY 0x00000008
#define RRF_RT_REG_DWORD 0x00000010
#define RRF_RT_REG_MULTI_SZ 0x00000020
#define RRF_RT_REG_QWORD 0x00000040
#define RRF_RT_DWORD (RRF_RT_REG_BINARY | RRF_RT_REG_DWORD)
#define RRF_RT_QWORD (RRF_RT_REG_BINARY | RRF_RT_REG_QWORD)
#define RRF_RT_ANY 0x0000ffff
#define RRF_NOEXPAND 0x10000000
#define RRF_ZEROONFAILURE 0x20000000
#define HKEY_CLASSES_ROOT PTR (_CAST,0x80000000)
#define HKEY_CURRENT_USER PTR (_CAST,0x80000001)
#define HKEY_LOCAL_MACHINE PTR (_CAST,0x80000002)
#define HKEY_USERS PTR (_CAST,0x80000003)
#define HKEY_PERFORMANCE_DATA PTR (_CAST,0x80000004)
#define HKEY_PERFORMANCE_TEXT PTR (_CAST,0x80000050)
#define HKEY_PERFORMANCE_NLSTEXT PTR (_CAST,0x80000060)
#define HKEY_CURRENT_CONFIG PTR (_CAST,0x80000005)
#define HKEY_DYN_DATA PTR (_CAST,0x80000006)
#define PROVIDER_KEEPS_VALUE_LENGTH 0x1
#define WIN31_CLASS NULL
#define FD_SETSIZE 64
#define IOCPARM_MASK 0x0000007f
#define IOC_VOID 0x20000000
#define IOC_OUT 0x40000000
#define IOC_IN 0x80000000
#define IOC_INOUT (IOC_IN|IOC_OUT)
#define IPPROTO_IP 0 
#define IPPROTO_HOPOPTS 0 
#define IPPROTO_ICMP 1 
#define IPPROTO_IGMP 2 
#define IPPROTO_GGP 3 
#define IPPROTO_IPV4 4 
#define IPPROTO_TCP 6 
#define IPPROTO_PUP 12 
#define IPPROTO_UDP 17 
#define IPPROTO_IDP 22 
#define IPPROTO_IPV6 41 
#define IPPROTO_ROUTING 43 
#define IPPROTO_FRAGMENT 44 
#define IPPROTO_ESP 50 
#define IPPROTO_AH 51 
#define IPPROTO_ICMPV6 58 
#define IPPROTO_NONE 59 
#define IPPROTO_DSTOPTS 60 
#define IPPROTO_ND 77 
#define IPPROTO_ICLFXBM 78
#define IPPROTO_RAW 255
#define IPPROTO_MAX 256
#define IPPORT_ECHO 7
#define IPPORT_DISCARD 9
#define IPPORT_SYSTAT 11
#define IPPORT_DAYTIME 13
#define IPPORT_NETSTAT 15
#define IPPORT_FTP 21
#define IPPORT_TELNET 23
#define IPPORT_SMTP 25
#define IPPORT_TIMESERVER 37
#define IPPORT_NAMESERVER 42
#define IPPORT_WHOIS 43
#define IPPORT_MTP 57
#define IPPORT_TFTP 69
#define IPPORT_RJE 77
#define IPPORT_FINGER 79
#define IPPORT_TTYLINK 87
#define IPPORT_SUPDUP 95
#define IPPORT_EXECSERVER 512
#define IPPORT_LOGINSERVER 513
#define IPPORT_CMDSERVER 514
#define IPPORT_EFSSERVER 520
#define IPPORT_BIFFUDP 512
#define IPPORT_WHOSERVER 513
#define IPPORT_ROUTESERVER 520
#define IPPORT_RESERVED 1024
#define IMPLINK_IP 155
#define IMPLINK_LOWEXPER 156
#define IMPLINK_HIGHEXPER 158
#define IN_CLASSA_NET 0xff000000
#define IN_CLASSA_NSHIFT 24
#define IN_CLASSA_HOST 0x00ffffff
#define IN_CLASSA_MAX 128
#define IN_CLASSB_NET 0xffff0000
#define IN_CLASSB_NSHIFT 16
#define IN_CLASSB_HOST 0x0000ffff
#define IN_CLASSB_MAX 65536
#define IN_CLASSC_NET 0xffffff00
#define IN_CLASSC_NSHIFT 8
#define IN_CLASSC_HOST 0x000000ff
#define INADDR_ANY DWORD(_CAST, 0x00000000)
#define INADDR_LOOPBACK 0x7f000001
#define INADDR_BROADCAST DWORD(_CAST, 0xffffffff)
#define INADDR_NONE 0xffffffff
#define WSADESCRIPTION_LEN 256
#define WSASYS_STATUS_LEN 128
#define IP_OPTIONS 1
#define IP_MULTICAST_IF 2
#define IP_MULTICAST_TTL 3
#define IP_MULTICAST_LOOP 4
#define IP_ADD_MEMBERSHIP 5
#define IP_DROP_MEMBERSHIP 6
#define IP_TTL 7 
#define IP_TOS 8 
#define IP_DONTFRAGMENT 9 
#define IP_DEFAULT_MULTICAST_TTL 1
#define IP_DEFAULT_MULTICAST_LOOP 1
#define IP_MAX_MEMBERSHIPS 20
#define INVALID_SOCKET DWORD(_CAST, 0xFFFFFFFF)
#define SOCKET_ERROR (-1)
#define FROM_PROTOCOL_INFO (-1)
#define SOCK_STREAM 1
#define SOCK_DGRAM 2
#define SOCK_RAW 3
#define SOCK_RDM 4
#define SOCK_SEQPACKET 5
#define SO_DEBUG 0x0001
#define SO_ACCEPTCONN 0x0002
#define SO_REUSEADDR 0x0004
#define SO_KEEPALIVE 0x0008
#define SO_DONTROUTE 0x0010
#define SO_BROADCAST 0x0020
#define SO_USELOOPBACK 0x0040
#define SO_LINGER 0x0080
#define SO_OOBINLINE 0x0100
#define SO_DONTLINGER DWORD(_CAST, 0xff7f)
#define SO_SNDBUF 0x1001
#define SO_RCVBUF 0x1002
#define SO_SNDLOWAT 0x1003
#define SO_RCVLOWAT 0x1004
#define SO_SNDTIMEO 0x1005
#define SO_RCVTIMEO 0x1006
#define SO_ERROR 0x1007
#define SO_TYPE 0x1008
#define SO_GROUP_ID 0x2001 
#define SO_GROUP_PRIORITY 0x2002 
#define SO_MAX_MSG_SIZE 0x2003 
#define SO_PROTOCOL_INFOA 0x2004 
#define SO_PROTOCOL_INFOW 0x2005 
#define SO_CONNDATA 0x7000
#define SO_CONNOPT 0x7001
#define SO_DISCDATA 0x7002
#define SO_DISCOPT 0x7003
#define SO_CONNDATALEN 0x7004
#define SO_CONNOPTLEN 0x7005
#define SO_DISCDATALEN 0x7006
#define SO_DISCOPTLEN 0x7007
#define SO_OPENTYPE 0x7008
#define SO_SYNCHRONOUS_ALERT 0x10
#define SO_SYNCHRONOUS_NONALERT 0x20
#define SO_MAXDG 0x7009
#define SO_MAXPATHDG 0x700A
#define SO_UPDATE_ACCEPT_CONTEXT 0x700B
#define SO_CONNECT_TIME 0x700C
#define TCP_NODELAY 0x0001
#define TCP_BSDURGENT 0x7000
#define AF_UNSPEC 0
#define AF_UNIX 1
#define AF_INET 2
#define AF_IMPLINK 3
#define AF_PUP 4
#define AF_CHAOS 5
#define AF_IPX 6
#define AF_NS 6
#define AF_ISO 7
#define AF_OSI AF_ISO
#define AF_ECMA 8
#define AF_DATAKIT 9
#define AF_CCITT 10
#define AF_SNA 11
#define AF_DECnet 12
#define AF_DLI 13
#define AF_LAT 14
#define AF_HYLINK 15
#define AF_APPLETALK 16
#define AF_NETBIOS 17
#define AF_VOICEVIEW 18
#define AF_FIREFOX 19 
#define AF_UNKNOWN1 20 
#define AF_BAN 21 
#define AF_ATM 22 
#define AF_INET6 23 
#define AF_CLUSTER 24 
#define AF_12844 25 
#define AF_IRDA 26 
#define AF_NETDES 28 
#define AF_TCNPROCESS 29
#define AF_TCNMESSAGE 30
#define AF_ICLFXBM 31
#define AF_MAX 32
#define _SS_MAXSIZE 128
#define PF_UNSPEC AF_UNSPEC
#define PF_UNIX AF_UNIX
#define PF_INET AF_INET
#define PF_IMPLINK AF_IMPLINK
#define PF_PUP AF_PUP
#define PF_CHAOS AF_CHAOS
#define PF_NS AF_NS
#define PF_IPX AF_IPX
#define PF_ISO AF_ISO
#define PF_OSI AF_OSI
#define PF_ECMA AF_ECMA
#define PF_DATAKIT AF_DATAKIT
#define PF_CCITT AF_CCITT
#define PF_SNA AF_SNA
#define PF_DECnet AF_DECnet
#define PF_DLI AF_DLI
#define PF_LAT AF_LAT
#define PF_HYLINK AF_HYLINK
#define PF_APPLETALK AF_APPLETALK
#define PF_VOICEVIEW AF_VOICEVIEW
#define PF_FIREFOX AF_FIREFOX
#define PF_UNKNOWN1 AF_UNKNOWN1
#define PF_BAN AF_BAN
#define PF_ATM AF_ATM
#define PF_INET6 AF_INET6
#define PF_MAX AF_MAX
#define SOL_SOCKET 0xffff
#define SOMAXCONN 0x7fffffff
#define MSG_OOB 0x1
#define MSG_PEEK 0x2
#define MSG_DONTROUTE 0x4
#define MSG_WAITALL 0x8 
#define MSG_PARTIAL 0x8000 
#define MSG_INTERRUPT 0x10 
#define MSG_MAXIOVLEN 16
#define MAXGETHOSTSTRUCT 1024
#define FD_READ_BIT 0
#define FD_READ (1 << FD_READ_BIT)
#define FD_WRITE_BIT 1
#define FD_WRITE (1 << FD_WRITE_BIT)
#define FD_OOB_BIT 2
#define FD_OOB (1 << FD_OOB_BIT)
#define FD_ACCEPT_BIT 3
#define FD_ACCEPT (1 << FD_ACCEPT_BIT)
#define FD_CONNECT_BIT 4
#define FD_CONNECT (1 << FD_CONNECT_BIT)
#define FD_CLOSE_BIT 5
#define FD_CLOSE (1 << FD_CLOSE_BIT)
#define FD_QOS_BIT 6
#define FD_QOS (1 << FD_QOS_BIT)
#define FD_GROUP_QOS_BIT 7
#define FD_GROUP_QOS (1 << FD_GROUP_QOS_BIT)
#define FD_ROUTING_INTERFACE_CHANGE_BIT 8
#define FD_ROUTING_INTERFACE_CHANGE (1 << FD_ROUTING_INTERFACE_CHANGE_BIT)
#define FD_ADDRESS_LIST_CHANGE_BIT 9
#define FD_ADDRESS_LIST_CHANGE (1 << FD_ADDRESS_LIST_CHANGE_BIT)
#define FD_MAX_EVENTS 10
#define FD_ALL_EVENTS ((1 << FD_MAX_EVENTS) - 1)
#define WSABASEERR 10000
#define WSAEINTR (WSABASEERR+4)
#define WSAEBADF (WSABASEERR+9)
#define WSAEACCES (WSABASEERR+13)
#define WSAEFAULT (WSABASEERR+14)
#define WSAEINVAL (WSABASEERR+22)
#define WSAEMFILE (WSABASEERR+24)
#define WSAEWOULDBLOCK (WSABASEERR+35)
#define WSAEINPROGRESS (WSABASEERR+36)
#define WSAEALREADY (WSABASEERR+37)
#define WSAENOTSOCK (WSABASEERR+38)
#define WSAEDESTADDRREQ (WSABASEERR+39)
#define WSAEMSGSIZE (WSABASEERR+40)
#define WSAEPROTOTYPE (WSABASEERR+41)
#define WSAENOPROTOOPT (WSABASEERR+42)
#define WSAEPROTONOSUPPORT (WSABASEERR+43)
#define WSAESOCKTNOSUPPORT (WSABASEERR+44)
#define WSAEOPNOTSUPP (WSABASEERR+45)
#define WSAEPFNOSUPPORT (WSABASEERR+46)
#define WSAEAFNOSUPPORT (WSABASEERR+47)
#define WSAEADDRINUSE (WSABASEERR+48)
#define WSAEADDRNOTAVAIL (WSABASEERR+49)
#define WSAENETDOWN (WSABASEERR+50)
#define WSAENETUNREACH (WSABASEERR+51)
#define WSAENETRESET (WSABASEERR+52)
#define WSAECONNABORTED (WSABASEERR+53)
#define WSAECONNRESET (WSABASEERR+54)
#define WSAENOBUFS (WSABASEERR+55)
#define WSAEISCONN (WSABASEERR+56)
#define WSAENOTCONN (WSABASEERR+57)
#define WSAESHUTDOWN (WSABASEERR+58)
#define WSAETOOMANYREFS (WSABASEERR+59)
#define WSAETIMEDOUT (WSABASEERR+60)
#define WSAECONNREFUSED (WSABASEERR+61)
#define WSAELOOP (WSABASEERR+62)
#define WSAENAMETOOLONG (WSABASEERR+63)
#define WSAEHOSTDOWN (WSABASEERR+64)
#define WSAEHOSTUNREACH (WSABASEERR+65)
#define WSAENOTEMPTY (WSABASEERR+66)
#define WSAEPROCLIM (WSABASEERR+67)
#define WSAEUSERS (WSABASEERR+68)
#define WSAEDQUOT (WSABASEERR+69)
#define WSAESTALE (WSABASEERR+70)
#define WSAEREMOTE (WSABASEERR+71)
#define WSASYSNOTREADY (WSABASEERR+91)
#define WSAVERNOTSUPPORTED (WSABASEERR+92)
#define WSANOTINITIALISED (WSABASEERR+93)
#define WSAEDISCON (WSABASEERR+101)
#define WSAENOMORE (WSABASEERR+102)
#define WSAECANCELLED (WSABASEERR+103)
#define WSAEINVALIDPROCTABLE (WSABASEERR+104)
#define WSAEINVALIDPROVIDER (WSABASEERR+105)
#define WSAEPROVIDERFAILEDINIT (WSABASEERR+106)
#define WSASYSCALLFAILURE (WSABASEERR+107)
#define WSASERVICE_NOT_FOUND (WSABASEERR+108)
#define WSATYPE_NOT_FOUND (WSABASEERR+109)
#define WSA_E_NO_MORE (WSABASEERR+110)
#define WSA_E_CANCELLED (WSABASEERR+111)
#define WSAEREFUSED (WSABASEERR+112)
#define WSAHOST_NOT_FOUND (WSABASEERR+1001)
#define HOST_NOT_FOUND WSAHOST_NOT_FOUND
#define WSATRY_AGAIN (WSABASEERR+1002)
#define WSANO_RECOVERY (WSABASEERR+1003)
#define WSANO_DATA (WSABASEERR+1004)
#define WSA_QOS_RECEIVERS (WSABASEERR + 1005)
#define WSA_QOS_SENDERS (WSABASEERR + 1006)
#define WSA_QOS_NO_SENDERS (WSABASEERR + 1007)
#define WSA_QOS_NO_RECEIVERS (WSABASEERR + 1008)
#define WSA_QOS_REQUEST_CONFIRMED (WSABASEERR + 1009)
#define WSA_QOS_ADMISSION_FAILURE (WSABASEERR + 1010)
#define WSA_QOS_POLICY_FAILURE (WSABASEERR + 1011)
#define WSA_QOS_BAD_STYLE (WSABASEERR + 1012)
#define WSA_QOS_BAD_OBJECT (WSABASEERR + 1013)
#define WSA_QOS_TRAFFIC_CTRL_ERROR (WSABASEERR + 1014)
#define WSA_QOS_GENERIC_ERROR (WSABASEERR + 1015)
#define WSA_QOS_ESERVICETYPE (WSABASEERR + 1016)
#define WSA_QOS_EFLOWSPEC (WSABASEERR + 1017)
#define WSA_QOS_EPROVSPECBUF (WSABASEERR + 1018)
#define WSA_QOS_EFILTERSTYLE (WSABASEERR + 1019)
#define WSA_QOS_EFILTERTYPE (WSABASEERR + 1020)
#define WSA_QOS_EFILTERCOUNT (WSABASEERR + 1021)
#define WSA_QOS_EOBJLENGTH (WSABASEERR + 1022)
#define WSA_QOS_EFLOWCOUNT (WSABASEERR + 1023)
#define WSA_QOS_EUNKOWNPSOBJ (WSABASEERR + 1024)
#define WSA_QOS_EPOLICYOBJ (WSABASEERR + 1025)
#define WSA_QOS_EFLOWDESC (WSABASEERR + 1026)
#define WSA_QOS_EPSFLOWSPEC (WSABASEERR + 1027)
#define WSA_QOS_EPSFILTERSPEC (WSABASEERR + 1028)
#define WSA_QOS_ESDMODEOBJ (WSABASEERR + 1029)
#define WSA_QOS_ESHAPERATEOBJ (WSABASEERR + 1030)
#define WSA_QOS_RESERVED_PETYPE (WSABASEERR + 1031)
#define TRY_AGAIN WSATRY_AGAIN
#define NO_RECOVERY WSANO_RECOVERY
#define NO_DATA WSANO_DATA
#define WSANO_ADDRESS WSANO_DATA
#define NO_ADDRESS WSANO_ADDRESS
#define CF_ACCEPT 0x0000
#define CF_REJECT 0x0001
#define CF_DEFER 0x0002
#define SD_RECEIVE 0x00
#define SD_SEND 0x01
#define SD_BOTH 0x02
#define SG_UNCONSTRAINED_GROUP 0x01
#define SG_CONSTRAINED_GROUP 0x02
#define MAX_PROTOCOL_CHAIN 7
#define BASE_PROTOCOL 1
#define LAYERED_PROTOCOL 0
#define JL_SENDER_ONLY 0x01
#define JL_RECEIVER_ONLY 0x02
#define JL_BOTH 0x04
#define WSA_FLAG_OVERLAPPED 0x01
#define WSA_FLAG_MULTIPOINT_C_ROOT 0x02
#define WSA_FLAG_MULTIPOINT_C_LEAF 0x04
#define WSA_FLAG_MULTIPOINT_D_ROOT 0x08
#define WSA_FLAG_MULTIPOINT_D_LEAF 0x10
#define IOC_UNIX 0x00000000
#define IOC_WS2 0x08000000
#define IOC_PROTOCOL 0x10000000
#define IOC_VENDOR 0x18000000
#define SERVICE_MULTIPLE (0x00000001)
#define NS_ALL (0)
#define NS_SAP (1)
#define NS_NDS (2)
#define NS_PEER_BROWSE (3)
#define NS_SLP (5)
#define NS_DHCP (6)
#define NS_TCPIP_LOCAL (10)
#define NS_TCPIP_HOSTS (11)
#define NS_DNS (12)
#define NS_NETBT (13)
#define NS_WINS (14)
#define NS_NLA (15) 
#define NS_NBP (20)
#define NS_MS (30)
#define NS_STDA (31)
#define NS_NTDS (32)
#define NS_X500 (40)
#define NS_NIS (41)
#define NS_NISPLUS (42)
#define NS_WRQ (50)
#define NS_NETDES (60) 
#define RES_UNUSED_1 (0x00000001)
#define RES_FLUSH_CACHE (0x00000002)
#define RES_SERVICE (0x00000004)
#define PRINTER_CONTROL_PAUSE 1
#define PRINTER_CONTROL_RESUME 2
#define PRINTER_CONTROL_PURGE 3
#define PRINTER_CONTROL_SET_STATUS 4
#define PRINTER_STATUS_PAUSED 0x00000001
#define PRINTER_STATUS_ERROR 0x00000002
#define PRINTER_STATUS_PENDING_DELETION 0x00000004
#define PRINTER_STATUS_PAPER_JAM 0x00000008
#define PRINTER_STATUS_PAPER_OUT 0x00000010
#define PRINTER_STATUS_MANUAL_FEED 0x00000020
#define PRINTER_STATUS_PAPER_PROBLEM 0x00000040
#define PRINTER_STATUS_OFFLINE 0x00000080
#define PRINTER_STATUS_IO_ACTIVE 0x00000100
#define PRINTER_STATUS_BUSY 0x00000200
#define PRINTER_STATUS_PRINTING 0x00000400
#define PRINTER_STATUS_OUTPUT_BIN_FULL 0x00000800
#define PRINTER_STATUS_NOT_AVAILABLE 0x00001000
#define PRINTER_STATUS_WAITING 0x00002000
#define PRINTER_STATUS_PROCESSING 0x00004000
#define PRINTER_STATUS_INITIALIZING 0x00008000
#define PRINTER_STATUS_WARMING_UP 0x00010000
#define PRINTER_STATUS_TONER_LOW 0x00020000
#define PRINTER_STATUS_NO_TONER 0x00040000
#define PRINTER_STATUS_PAGE_PUNT 0x00080000
#define PRINTER_STATUS_USER_INTERVENTION 0x00100000
#define PRINTER_STATUS_OUT_OF_MEMORY 0x00200000
#define PRINTER_STATUS_DOOR_OPEN 0x00400000
#define PRINTER_STATUS_SERVER_UNKNOWN 0x00800000
#define PRINTER_STATUS_POWER_SAVE 0x01000000
#define PRINTER_ATTRIBUTE_QUEUED 0x00000001
#define PRINTER_ATTRIBUTE_DIRECT 0x00000002
#define PRINTER_ATTRIBUTE_DEFAULT 0x00000004
#define PRINTER_ATTRIBUTE_SHARED 0x00000008
#define PRINTER_ATTRIBUTE_NETWORK 0x00000010
#define PRINTER_ATTRIBUTE_HIDDEN 0x00000020
#define PRINTER_ATTRIBUTE_LOCAL 0x00000040
#define PRINTER_ATTRIBUTE_ENABLE_DEVQ 0x00000080
#define PRINTER_ATTRIBUTE_KEEPPRINTEDJOBS 0x00000100
#define PRINTER_ATTRIBUTE_DO_COMPLETE_FIRST 0x00000200
#define PRINTER_ATTRIBUTE_WORK_OFFLINE 0x00000400
#define PRINTER_ATTRIBUTE_ENABLE_BIDI 0x00000800
#define PRINTER_ATTRIBUTE_RAW_ONLY 0x00001000
#define PRINTER_ATTRIBUTE_PUBLISHED 0x00002000
#define PRINTER_ATTRIBUTE_FAX 0x00004000
#define PRINTER_ATTRIBUTE_TS 0x00008000
#define NO_PRIORITY 0
#define MAX_PRIORITY 99
#define MIN_PRIORITY 1
#define DEF_PRIORITY 1
#define JOB_CONTROL_PAUSE 1
#define JOB_CONTROL_RESUME 2
#define JOB_CONTROL_CANCEL 3
#define JOB_CONTROL_RESTART 4
#define JOB_CONTROL_DELETE 5
#define JOB_CONTROL_SENT_TO_PRINTER 6
#define JOB_CONTROL_LAST_PAGE_EJECTED 7
#define JOB_STATUS_PAUSED 0x00000001
#define JOB_STATUS_ERROR 0x00000002
#define JOB_STATUS_DELETING 0x00000004
#define JOB_STATUS_SPOOLING 0x00000008
#define JOB_STATUS_PRINTING 0x00000010
#define JOB_STATUS_OFFLINE 0x00000020
#define JOB_STATUS_PAPEROUT 0x00000040
#define JOB_STATUS_PRINTED 0x00000080
#define JOB_STATUS_DELETED 0x00000100
#define JOB_STATUS_BLOCKED_DEVQ 0x00000200
#define JOB_STATUS_USER_INTERVENTION 0x00000400
#define JOB_STATUS_RESTART 0x00000800
#define JOB_STATUS_COMPLETE 0x00001000
#define JOB_POSITION_UNSPECIFIED 0
#define DI_CHANNEL 1
#define DI_CHANNEL_WRITE 2
#define DI_READ_SPOOL_JOB 3
#define FORM_BUILTIN 0x00000001
#define PORT_TYPE_WRITE 0x0001
#define PORT_TYPE_READ 0x0002
#define PORT_TYPE_REDIRECTED 0x0004
#define PORT_TYPE_NET_ATTACHED 0x0008
#define PORT_STATUS_TYPE_ERROR 1
#define PORT_STATUS_TYPE_WARNING 2
#define PORT_STATUS_TYPE_INFO 3
#define PORT_STATUS_OFFLINE 1
#define PORT_STATUS_PAPER_JAM 2
#define PORT_STATUS_PAPER_OUT 3
#define PORT_STATUS_OUTPUT_BIN_FULL 4
#define PORT_STATUS_PAPER_PROBLEM 5
#define PORT_STATUS_NO_TONER 6
#define PORT_STATUS_DOOR_OPEN 7
#define PORT_STATUS_USER_INTERVENTION 8
#define PORT_STATUS_OUT_OF_MEMORY 9
#define PORT_STATUS_TONER_LOW 10
#define PORT_STATUS_WARMING_UP 11
#define PORT_STATUS_POWER_SAVE 12
#define PRINTER_ENUM_DEFAULT 0x00000001
#define PRINTER_ENUM_LOCAL 0x00000002
#define PRINTER_ENUM_CONNECTIONS 0x00000004
#define PRINTER_ENUM_FAVORITE 0x00000004
#define PRINTER_ENUM_NAME 0x00000008
#define PRINTER_ENUM_REMOTE 0x00000010
#define PRINTER_ENUM_SHARED 0x00000020
#define PRINTER_ENUM_NETWORK 0x00000040
#define PRINTER_ENUM_EXPAND 0x00004000
#define PRINTER_ENUM_CONTAINER 0x00008000
#define PRINTER_ENUM_ICONMASK 0x00ff0000
#define PRINTER_ENUM_ICON1 0x00010000
#define PRINTER_ENUM_ICON2 0x00020000
#define PRINTER_ENUM_ICON3 0x00040000
#define PRINTER_ENUM_ICON4 0x00080000
#define PRINTER_ENUM_ICON5 0x00100000
#define PRINTER_ENUM_ICON6 0x00200000
#define PRINTER_ENUM_ICON7 0x00400000
#define PRINTER_ENUM_ICON8 0x00800000
#define PRINTER_ENUM_HIDE 0x01000000
#define SPOOL_FILE_PERSISTENT 0x00000001
#define SPOOL_FILE_TEMPORARY 0x00000002
#define PRINTER_NOTIFY_TYPE 0x00
#define JOB_NOTIFY_TYPE 0x01
#define PRINTER_NOTIFY_FIELD_SERVER_NAME 0x00
#define PRINTER_NOTIFY_FIELD_PRINTER_NAME 0x01
#define PRINTER_NOTIFY_FIELD_SHARE_NAME 0x02
#define PRINTER_NOTIFY_FIELD_PORT_NAME 0x03
#define PRINTER_NOTIFY_FIELD_DRIVER_NAME 0x04
#define PRINTER_NOTIFY_FIELD_COMMENT 0x05
#define PRINTER_NOTIFY_FIELD_LOCATION 0x06
#define PRINTER_NOTIFY_FIELD_DEVMODE 0x07
#define PRINTER_NOTIFY_FIELD_SEPFILE 0x08
#define PRINTER_NOTIFY_FIELD_PRINT_PROCESSOR 0x09
#define PRINTER_NOTIFY_FIELD_PARAMETERS 0x0A
#define PRINTER_NOTIFY_FIELD_DATATYPE 0x0B
#define PRINTER_NOTIFY_FIELD_SECURITY_DESCRIPTOR 0x0C
#define PRINTER_NOTIFY_FIELD_ATTRIBUTES 0x0D
#define PRINTER_NOTIFY_FIELD_PRIORITY 0x0E
#define PRINTER_NOTIFY_FIELD_DEFAULT_PRIORITY 0x0F
#define PRINTER_NOTIFY_FIELD_START_TIME 0x10
#define PRINTER_NOTIFY_FIELD_UNTIL_TIME 0x11
#define PRINTER_NOTIFY_FIELD_STATUS 0x12
#define PRINTER_NOTIFY_FIELD_STATUS_STRING 0x13
#define PRINTER_NOTIFY_FIELD_CJOBS 0x14
#define PRINTER_NOTIFY_FIELD_AVERAGE_PPM 0x15
#define PRINTER_NOTIFY_FIELD_TOTAL_PAGES 0x16
#define PRINTER_NOTIFY_FIELD_PAGES_PRINTED 0x17
#define PRINTER_NOTIFY_FIELD_TOTAL_BYTES 0x18
#define PRINTER_NOTIFY_FIELD_BYTES_PRINTED 0x19
#define PRINTER_NOTIFY_FIELD_OBJECT_GUID 0x1A
#define JOB_NOTIFY_FIELD_PRINTER_NAME 0x00
#define JOB_NOTIFY_FIELD_MACHINE_NAME 0x01
#define JOB_NOTIFY_FIELD_PORT_NAME 0x02
#define JOB_NOTIFY_FIELD_USER_NAME 0x03
#define JOB_NOTIFY_FIELD_NOTIFY_NAME 0x04
#define JOB_NOTIFY_FIELD_DATATYPE 0x05
#define JOB_NOTIFY_FIELD_PRINT_PROCESSOR 0x06
#define JOB_NOTIFY_FIELD_PARAMETERS 0x07
#define JOB_NOTIFY_FIELD_DRIVER_NAME 0x08
#define JOB_NOTIFY_FIELD_DEVMODE 0x09
#define JOB_NOTIFY_FIELD_STATUS 0x0A
#define JOB_NOTIFY_FIELD_STATUS_STRING 0x0B
#define JOB_NOTIFY_FIELD_SECURITY_DESCRIPTOR 0x0C
#define JOB_NOTIFY_FIELD_DOCUMENT 0x0D
#define JOB_NOTIFY_FIELD_PRIORITY 0x0E
#define JOB_NOTIFY_FIELD_POSITION 0x0F
#define JOB_NOTIFY_FIELD_SUBMITTED 0x10
#define JOB_NOTIFY_FIELD_START_TIME 0x11
#define JOB_NOTIFY_FIELD_UNTIL_TIME 0x12
#define JOB_NOTIFY_FIELD_TIME 0x13
#define JOB_NOTIFY_FIELD_TOTAL_PAGES 0x14
#define JOB_NOTIFY_FIELD_PAGES_PRINTED 0x15
#define JOB_NOTIFY_FIELD_TOTAL_BYTES 0x16
#define JOB_NOTIFY_FIELD_BYTES_PRINTED 0x17
#define PRINTER_NOTIFY_OPTIONS_REFRESH 0x01
#define PRINTER_NOTIFY_INFO_DISCARDED 0x01
#define PRINTER_CHANGE_ADD_PRINTER 0x00000001
#define PRINTER_CHANGE_SET_PRINTER 0x00000002
#define PRINTER_CHANGE_DELETE_PRINTER 0x00000004
#define PRINTER_CHANGE_FAILED_CONNECTION_PRINTER 0x00000008
#define PRINTER_CHANGE_PRINTER 0x000000FF
#define PRINTER_CHANGE_ADD_JOB 0x00000100
#define PRINTER_CHANGE_SET_JOB 0x00000200
#define PRINTER_CHANGE_DELETE_JOB 0x00000400
#define PRINTER_CHANGE_WRITE_JOB 0x00000800
#define PRINTER_CHANGE_JOB 0x0000FF00
#define PRINTER_CHANGE_ADD_FORM 0x00010000
#define PRINTER_CHANGE_SET_FORM 0x00020000
#define PRINTER_CHANGE_DELETE_FORM 0x00040000
#define PRINTER_CHANGE_FORM 0x00070000
#define PRINTER_CHANGE_ADD_PORT 0x00100000
#define PRINTER_CHANGE_CONFIGURE_PORT 0x00200000
#define PRINTER_CHANGE_DELETE_PORT 0x00400000
#define PRINTER_CHANGE_PORT 0x00700000
#define PRINTER_CHANGE_ADD_PRINT_PROCESSOR 0x01000000
#define PRINTER_CHANGE_DELETE_PRINT_PROCESSOR 0x04000000
#define PRINTER_CHANGE_PRINT_PROCESSOR 0x07000000
#define PRINTER_CHANGE_ADD_PRINTER_DRIVER 0x10000000
#define PRINTER_CHANGE_SET_PRINTER_DRIVER 0x20000000
#define PRINTER_CHANGE_DELETE_PRINTER_DRIVER 0x40000000
#define PRINTER_CHANGE_PRINTER_DRIVER 0x70000000
#define PRINTER_CHANGE_TIMEOUT 0x80000000
#define PRINTER_CHANGE_ALL 0x7777FFFF
#define PRINTER_ERROR_INFORMATION 0x80000000
#define PRINTER_ERROR_WARNING 0x40000000
#define PRINTER_ERROR_SEVERE 0x20000000
#define PRINTER_ERROR_OUTOFPAPER 0x00000001
#define PRINTER_ERROR_JAM 0x00000002
#define PRINTER_ERROR_OUTOFTONER 0x00000004
#define SERVER_ACCESS_ADMINISTER 0x00000001
#define SERVER_ACCESS_ENUMERATE 0x00000002
#define PRINTER_ACCESS_ADMINISTER 0x00000004
#define PRINTER_ACCESS_USE 0x00000008
#define JOB_ACCESS_ADMINISTER 0x00000010
#define JOB_ACCESS_READ 0x00000020
#define SERVER_ALL_ACCESS 0x000f0003
#define SERVER_READ 0x00020002
#define SERVER_WRITE 0x00020003
#define SERVER_EXECUTE 0x00020002
#define PRINTER_ALL_ACCESS 0x000f000c
#define PRINTER_READ 0x00020008
#define PRINTER_WRITE 0x00020008
#define PRINTER_EXECUTE 0x00020008
#define JOB_ALL_ACCESS 0x000f0010
#define JOB_READ 0x00020010
#define JOB_WRITE 0x00020010
#define JOB_EXECUTE 0x00020010
#define SERVICE_CONTROL_RUN 0x00000000
#define SERVICE_NO_CHANGE 0xFFFFFFFF
#define SERVICE_ACTIVE 0x00000001
#define SERVICE_INACTIVE 0x00000002
#define SERVICE_STATE_ALL 0x00000003
#define SERVICE_CONTROL_STOP 0x00000001
#define SERVICE_CONTROL_PAUSE 0x00000002
#define SERVICE_CONTROL_CONTINUE 0x00000003
#define SERVICE_CONTROL_INTERROGATE 0x00000004
#define SERVICE_CONTROL_SHUTDOWN 0x00000005
#define SERVICE_CONTROL_PARAMCHANGE 0x00000006
#define SERVICE_CONTROL_NETBINDADD 0x00000007
#define SERVICE_CONTROL_NETBINDREMOVE 0x00000008
#define SERVICE_CONTROL_NETBINDENABLE 0x00000009
#define SERVICE_CONTROL_NETBINDDISABLE 0x0000000A
#define SERVICE_CONTROL_DEVICEEVENT 0x0000000B
#define SERVICE_CONTROL_HARDWAREPROFILECHANGE 0x0000000C
#define SERVICE_CONTROL_POWEREVENT 0x0000000D
#define SERVICE_CONTROL_SESSIONCHANGE 0x0000000E
#define SERVICE_STOPPED 0x00000001
#define SERVICE_START_PENDING 0x00000002
#define SERVICE_STOP_PENDING 0x00000003
#define SERVICE_RUNNING 0x00000004
#define SERVICE_CONTINUE_PENDING 0x00000005
#define SERVICE_PAUSE_PENDING 0x00000006
#define SERVICE_PAUSED 0x00000007
#define SERVICE_ACCEPT_STOP 0x00000001
#define SERVICE_ACCEPT_PAUSE_CONTINUE 0x00000002
#define SERVICE_ACCEPT_SHUTDOWN 0x00000004
#define SERVICE_ACCEPT_PARAMCHANGE 0x00000008
#define SERVICE_ACCEPT_NETBINDCHANGE 0x00000010
#define SERVICE_ACCEPT_HARDWAREPROFILECHANGE 0x00000020
#define SERVICE_ACCEPT_POWEREVENT 0x00000040
#define SERVICE_ACCEPT_SESSIONCHANGE 0x00000080
#define SC_MANAGER_CONNECT 0x0001
#define SC_MANAGER_CREATE_SERVICE 0x0002
#define SC_MANAGER_ENUMERATE_SERVICE 0x0004
#define SC_MANAGER_LOCK 0x0008
#define SC_MANAGER_QUERY_LOCK_STATUS 0x0010
#define SC_MANAGER_MODIFY_BOOT_CONFIG 0x0020
#define SC_MANAGER_ALL_ACCESS 0x000F003FL
#define SERVICE_QUERY_CONFIG 0x0001
#define SERVICE_CHANGE_CONFIG 0x0002
#define SERVICE_QUERY_STATUS 0x0004
#define SERVICE_ENUMERATE_DEPENDENTS 0x0008
#define SERVICE_START 0x0010
#define SERVICE_STOP 0x0020
#define SERVICE_PAUSE_CONTINUE 0x0040
#define SERVICE_INTERROGATE 0x0080
#define SERVICE_USER_DEFINED_CONTROL 0x0100
#define SERVICE_ALL_ACCESS 0x000F01FFL
#define RC_RT_CURSOR 1
#define RC_RT_BITMAP 2
#define RC_RT_ICON 3
#define RC_RT_MENU 4
#define RC_RT_DIALOG 5
#define RC_RT_STRING 6
#define RC_RT_FONTDIR 7
#define RC_RT_FONT 8
#define RC_RT_ACCELERATOR 9
#define RC_RT_RCDATA 10
#define RC_RT_MESSAGETABLE 11
#define RC_RT_GROUP_CURSOR 12
#define RC_RT_GROUP_ICON 14
#define RC_RT_VERSION 16
#define RC_RT_DLGINCLUDE 17
#define RC_RT_PLUGPLAY 19
#define RC_RT_VXD 20
#define RC_RT_ANICURSOR 21
#define RC_RT_ANIICON 22
#define RC_RT_HTML 23
#define RC_RT_MANIFEST 24
#define RT_CURSOR PTR (_CAST,1)
#define RT_BITMAP PTR (_CAST,2)
#define RT_ICON PTR (_CAST,3)
#define RT_MENU PTR (_CAST,4)
#define RT_DIALOG PTR (_CAST,5)
#define RT_STRING PTR (_CAST,6)
#define RT_FONTDIR PTR (_CAST,7)
#define RT_FONT PTR (_CAST,8)
#define RT_ACCELERATOR PTR (_CAST,9)
#define RT_RCDATA PTR (_CAST,10)
#define RT_MESSAGETABLE PTR (_CAST,11)
#define DIFFERENCE 11
#define RT_GROUP_CURSOR PTR(_CAST, 12)
#define RT_GROUP_ICON PTR(_CAST, 14)
#define RT_VERSION PTR (_CAST,16)
#define RT_DLGINCLUDE PTR (_CAST,17)
#define RT_PLUGPLAY PTR (_CAST,19)
#define RT_VXD PTR (_CAST,20)
#define RT_ANICURSOR PTR (_CAST,21)
#define RT_ANIICON PTR (_CAST,22)
#define RT_HTML PTR (_CAST,23)
#define RT_MANIFEST PTR (_CAST,24)
#define CREATEPROCESS_MANIFEST_RESOURCE_ID 1
#define ISOLATIONAWARE_MANIFEST_RESOURCE_ID 2
#define ISOLATIONAWARE_NOSTATICIMPORT_MANIFEST_RESOURCE_ID 3
#define SB_HORZ 0
#define SB_VERT 1
#define SB_CTL 2
#define SB_BOTH 3
#define SB_LINEUP 0
#define SB_LINELEFT 0
#define SB_LINEDOWN 1
#define SB_LINERIGHT 1
#define SB_PAGEUP 2
#define SB_PAGELEFT 2
#define SB_PAGEDOWN 3
#define SB_PAGERIGHT 3
#define SB_THUMBPOSITION 4
#define SB_THUMBTRACK 5
#define SB_TOP 6
#define SB_LEFT 6
#define SB_BOTTOM 7
#define SB_RIGHT 7
#define SB_ENDSCROLL 8
#define SW_HIDE 0
#define SW_SHOWNORMAL 1
#define SW_NORMAL 1
#define SW_SHOWMINIMIZED 2
#define SW_SHOWMAXIMIZED 3
#define SW_MAXIMIZE 3
#define SW_SHOWNOACTIVATE 4
#define SW_SHOW 5
#define SW_MINIMIZE 6
#define SW_SHOWMINNOACTIVE 7
#define SW_SHOWNA 8
#define SW_RESTORE 9
#define SW_SHOWDEFAULT 10
#define SW_FORCEMINIMIZE 11
#define SW_MAX 11
#define HIDE_WINDOW 0
#define SHOW_OPENWINDOW 1
#define SHOW_ICONWINDOW 2
#define SHOW_FULLSCREEN 3
#define SHOW_OPENNOACTIVATE 4
#define SW_PARENTCLOSING 1
#define SW_OTHERZOOM 2
#define SW_PARENTOPENING 3
#define SW_OTHERUNZOOM 4
#define AW_HOR_POSITIVE 0x00000001
#define AW_HOR_NEGATIVE 0x00000002
#define AW_VER_POSITIVE 0x00000004
#define AW_VER_NEGATIVE 0x00000008
#define AW_CENTER 0x00000010
#define AW_HIDE 0x00010000
#define AW_ACTIVATE 0x00020000
#define AW_SLIDE 0x00040000
#define AW_BLEND 0x00080000
#define KF_EXTENDED 0x0100
#define KF_DLGMODE 0x0800
#define KF_MENUMODE 0x1000
#define KF_ALTDOWN 0x2000
#define KF_REPEAT 0x4000
#define KF_UP 0x8000
#define VK_LBUTTON 0x01
#define VK_RBUTTON 0x02
#define VK_CANCEL 0x03
#define VK_MBUTTON 0x04 
#define VK_XBUTTON1 0x05 
#define VK_XBUTTON2 0x06 
#define VK_BACK 0x08
#define VK_TAB 0x09
#define VK_CLEAR 0x0C
#define VK_RETURN 0x0D
#define VK_SHIFT 0x10
#define VK_CONTROL 0x11
#define VK_MENU 0x12
#define VK_PAUSE 0x13
#define VK_CAPITAL 0x14
#define VK_KANA 0x15
#define VK_HANGEUL 0x15 
#define VK_HANGUL 0x15
#define VK_JUNJA 0x17
#define VK_FINAL 0x18
#define VK_HANJA 0x19
#define VK_KANJI 0x19
#define VK_ESCAPE 0x1B
#define VK_CONVERT 0x1C
#define VK_NONCONVERT 0x1D
#define VK_ACCEPT 0x1E
#define VK_MODECHANGE 0x1F
#define VK_SPACE 0x20
#define VK_PRIOR 0x21
#define VK_NEXT 0x22
#define VK_END 0x23
#define VK_HOME 0x24
#define VK_LEFT 0x25
#define VK_UP 0x26
#define VK_RIGHT 0x27
#define VK_DOWN 0x28
#define VK_SELECT 0x29
#define VK_PRINT 0x2A
#define VK_EXECUTE 0x2B
#define VK_SNAPSHOT 0x2C
#define VK_INSERT 0x2D
#define VK_DELETE 0x2E
#define VK_HELP 0x2F
#define VK_LWIN 0x5B
#define VK_RWIN 0x5C
#define VK_APPS 0x5D
#define VK_SLEEP 0x5F
#define VK_NUMPAD0 0x60
#define VK_NUMPAD1 0x61
#define VK_NUMPAD2 0x62
#define VK_NUMPAD3 0x63
#define VK_NUMPAD4 0x64
#define VK_NUMPAD5 0x65
#define VK_NUMPAD6 0x66
#define VK_NUMPAD7 0x67
#define VK_NUMPAD8 0x68
#define VK_NUMPAD9 0x69
#define VK_MULTIPLY 0x6A
#define VK_ADD 0x6B
#define VK_SEPARATOR 0x6C
#define VK_SUBTRACT 0x6D
#define VK_DECIMAL 0x6E
#define VK_DIVIDE 0x6F
#define VK_F1 0x70
#define VK_F2 0x71
#define VK_F3 0x72
#define VK_F4 0x73
#define VK_F5 0x74
#define VK_F6 0x75
#define VK_F7 0x76
#define VK_F8 0x77
#define VK_F9 0x78
#define VK_F10 0x79
#define VK_F11 0x7A
#define VK_F12 0x7B
#define VK_F13 0x7C
#define VK_F14 0x7D
#define VK_F15 0x7E
#define VK_F16 0x7F
#define VK_F17 0x80
#define VK_F18 0x81
#define VK_F19 0x82
#define VK_F20 0x83
#define VK_F21 0x84
#define VK_F22 0x85
#define VK_F23 0x86
#define VK_F24 0x87
#define VK_NUMLOCK 0x90
#define VK_SCROLL 0x91
#define VK_OEM_SCROLL 0x91
#define VK_OEM_NEC_EQUAL 0x92
#define VK_OEM_FJ_JISHO 0x92
#define VK_OEM_FJ_MASSHOU 0x93
#define VK_OEM_FJ_TOUROKU 0x94
#define VK_OEM_FJ_LOYA 0x95
#define VK_OEM_FJ_ROYA 0x96
#define VK_LSHIFT 0xA0
#define VK_RSHIFT 0xA1
#define VK_LCONTROL 0xA2
#define VK_RCONTROL 0xA3
#define VK_LMENU 0xA4
#define VK_RMENU 0xA5
#define VK_BROWSER_BACK 0xA6
#define VK_BROWSER_FORWARD 0xA7
#define VK_BROWSER_REFRESH 0xA8
#define VK_BROWSER_STOP 0xA9
#define VK_BROWSER_SEARCH 0xAA
#define VK_BROWSER_FAVORITES 0xAB
#define VK_BROWSER_HOME 0xAC
#define VK_VOLUME_MUTE 0xAD
#define VK_VOLUME_DOWN 0xAE
#define VK_VOLUME_UP 0xAF
#define VK_MEDIA_NEXT_TRACK 0xB0
#define VK_MEDIA_PREV_TRACK 0xB1
#define VK_MEDIA_STOP 0xB2
#define VK_MEDIA_PLAY_PAUSE 0xB3
#define VK_LAUNCH_MAIL 0xB4
#define VK_LAUNCH_MEDIA_SELECT 0xB5
#define VK_LAUNCH_APP1 0xB6
#define VK_LAUNCH_APP2 0xB7
#define VK_OEM_1 0xBA
#define VK_OEM_PLUS 0xBB
#define VK_OEM_COMMA 0xBC
#define VK_OEM_MINUS 0xBD
#define VK_OEM_PERIOD 0xBE
#define VK_OEM_2 0xBF
#define VK_OEM_3 0xC0
#define VK_OEM_4 0xDB
#define VK_OEM_5 0xDC
#define VK_OEM_6 0xDD
#define VK_OEM_7 0xDE
#define VK_OEM_8 0xDF
#define VK_OEM_AX 0xE1
#define VK_OEM_102 0xE2
#define VK_ICO_HELP 0xE3
#define VK_ICO_00 0xE4
#define VK_PROCESSKEY 0xE5
#define VK_ICO_CLEAR 0xE6
#define VK_PACKET 0xE7
#define VK_OEM_RESET 0xE9
#define VK_OEM_JUMP 0xEA
#define VK_OEM_PA1 0xEB
#define VK_OEM_PA2 0xEC
#define VK_OEM_PA3 0xED
#define VK_OEM_WSCTRL 0xEE
#define VK_OEM_CUSEL 0xEF
#define VK_OEM_ATTN 0xF0
#define VK_OEM_FINISH 0xF1
#define VK_OEM_COPY 0xF2
#define VK_OEM_AUTO 0xF3
#define VK_OEM_ENLW 0xF4
#define VK_OEM_BACKTAB 0xF5
#define VK_ATTN 0xF6
#define VK_CRSEL 0xF7
#define VK_EXSEL 0xF8
#define VK_EREOF 0xF9
#define VK_PLAY 0xFA
#define VK_ZOOM 0xFB
#define VK_NONAME 0xFC
#define VK_PA1 0xFD
#define VK_OEM_CLEAR 0xFE
#define WH_MIN (-1)
#define WH_MSGFILTER (-1)
#define WH_JOURNALRECORD 0
#define WH_JOURNALPLAYBACK 1
#define WH_KEYBOARD 2
#define WH_GETMESSAGE 3
#define WH_CALLWNDPROC 4
#define WH_CBT 5
#define WH_SYSMSGFILTER 6
#define WH_MOUSE 7
#define WH_HARDWARE 8
#define WH_DEBUG 9
#define WH_SHELL 10
#define WH_FOREGROUNDIDLE 11
#define WH_CALLWNDPROCRET 12
#define WH_KEYBOARD_LL 13
#define WH_MOUSE_LL 14
#define WH_MAX 14
#define WH_MINHOOK WH_MIN
#define WH_MAXHOOK WH_MAX
#define HC_ACTION 0
#define HC_GETNEXT 1
#define HC_SKIP 2
#define HC_NOREMOVE 3
#define HC_NOREM HC_NOREMOVE
#define HC_SYSMODALON 4
#define HC_SYSMODALOFF 5
#define HCBT_MOVESIZE 0
#define HCBT_MINMAX 1
#define HCBT_QS 2
#define HCBT_CREATEWND 3
#define HCBT_DESTROYWND 4
#define HCBT_ACTIVATE 5
#define HCBT_CLICKSKIPPED 6
#define HCBT_KEYSKIPPED 7
#define HCBT_SYSCOMMAND 8
#define HCBT_SETFOCUS 9
#define MSGF_DIALOGBOX 0
#define MSGF_MESSAGEBOX 1
#define MSGF_MENU 2
#define MSGF_MOVE 3
#define MSGF_SIZE 4
#define MSGF_SCROLLBAR 5
#define MSGF_NEXTWINDOW 6
#define MSGF_MAINLOOP 8
#define MSGF_MAX 8
#define MSGF_USER 4096
#define HSHELL_WINDOWCREATED 1
#define HSHELL_WINDOWDESTROYED 2
#define HSHELL_ACTIVATESHELLWINDOW 3
#define HSHELL_WINDOWACTIVATED 4
#define HSHELL_GETMINRECT 5
#define HSHELL_REDRAW 6
#define HSHELL_TASKMAN 7
#define HSHELL_LANGUAGE 8
#define HSHELL_SYSMENU 9
#define HSHELL_ENDTASK 10
#define HSHELL_ACCESSIBILITYSTATE 11
#define HSHELL_APPCOMMAND 12
#define HSHELL_WINDOWREPLACED 13
#define HSHELL_WINDOWREPLACING 14
#define HSHELL_HIGHBIT 0x8000
#define HSHELL_FLASH 0x8005
#define HSHELL_RUDEAPPACTIVATED 0x8004
#define ACCESS_STICKYKEYS 0x0001
#define ACCESS_FILTERKEYS 0x0002
#define ACCESS_MOUSEKEYS 0x0003
#define APPCOMMAND_BROWSER_BACKWARD 1
#define APPCOMMAND_BROWSER_FORWARD 2
#define APPCOMMAND_BROWSER_REFRESH 3
#define APPCOMMAND_BROWSER_STOP 4
#define APPCOMMAND_BROWSER_SEARCH 5
#define APPCOMMAND_BROWSER_FAVORITES 6
#define APPCOMMAND_BROWSER_HOME 7
#define APPCOMMAND_VOLUME_MUTE 8
#define APPCOMMAND_VOLUME_DOWN 9
#define APPCOMMAND_VOLUME_UP 10
#define APPCOMMAND_MEDIA_NEXTTRACK 11
#define APPCOMMAND_MEDIA_PREVIOUSTRACK 12
#define APPCOMMAND_MEDIA_STOP 13
#define APPCOMMAND_MEDIA_PLAY_PAUSE 14
#define APPCOMMAND_LAUNCH_MAIL 15
#define APPCOMMAND_LAUNCH_MEDIA_SELECT 16
#define APPCOMMAND_LAUNCH_APP1 17
#define APPCOMMAND_LAUNCH_APP2 18
#define APPCOMMAND_BASS_DOWN 19
#define APPCOMMAND_BASS_BOOST 20
#define APPCOMMAND_BASS_UP 21
#define APPCOMMAND_TREBLE_DOWN 22
#define APPCOMMAND_TREBLE_UP 23
#define APPCOMMAND_MICROPHONE_VOLUME_MUTE 24
#define APPCOMMAND_MICROPHONE_VOLUME_DOWN 25
#define APPCOMMAND_MICROPHONE_VOLUME_UP 26
#define APPCOMMAND_HELP 27
#define APPCOMMAND_FIND 28
#define APPCOMMAND_NEW 29
#define APPCOMMAND_OPEN 30
#define APPCOMMAND_CLOSE 31
#define APPCOMMAND_SAVE 32
#define APPCOMMAND_PRINT 33
#define APPCOMMAND_UNDO 34
#define APPCOMMAND_REDO 35
#define APPCOMMAND_COPY 36
#define APPCOMMAND_CUT 37
#define APPCOMMAND_PASTE 38
#define APPCOMMAND_REPLY_TO_MAIL 39
#define APPCOMMAND_FORWARD_MAIL 40
#define APPCOMMAND_SEND_MAIL 41
#define APPCOMMAND_SPELL_CHECK 42
#define APPCOMMAND_DICTATE_OR_COMMAND_CONTROL_TOGGLE 43
#define APPCOMMAND_MIC_ON_OFF_TOGGLE 44
#define APPCOMMAND_CORRECTION_LIST 45
#define APPCOMMAND_MEDIA_CHANNEL_DOWN 52
#define APPCOMMAND_MEDIA_CHANNEL_UP 51
#define APPCOMMAND_MEDIA_FASTFORWARD 49
#define APPCOMMAND_MEDIA_PAUSE 47
#define APPCOMMAND_MEDIA_PLAY 46
#define APPCOMMAND_MEDIA_RECORD 48
#define APPCOMMAND_MEDIA_REWIND 50
#define FAPPCOMMAND_KEY 0
#define FAPPCOMMAND_MOUSE 0x8000
#define FAPPCOMMAND_OEM 0x1000
#define FAPPCOMMAND_MASK 0xF000
#define HKL_PREV 0
#define HKL_NEXT 1
#define KLF_ACTIVATE 0x00000001
#define KLF_SUBSTITUTE_OK 0x00000002
#define KLF_UNLOADPREVIOUS 0x00000004
#define KLF_REORDER 0x00000008
#define KLF_REPLACELANG 0x00000010
#define KLF_NOTELLSHELL 0x00000080
#define KLF_SETFORPROCESS 0x00000100
#define KLF_SHIFTLOCK 0x00010000
#define KLF_RESET 0x40000000
#define KL_NAMELENGTH 9
#define DESKTOP_READOBJECTS 0x0001L
#define DESKTOP_CREATEWINDOW 0x0002L
#define DESKTOP_CREATEMENU 0x0004L
#define DESKTOP_HOOKCONTROL 0x0008L
#define DESKTOP_JOURNALRECORD 0x0010L
#define DESKTOP_JOURNALPLAYBACK 0x0020L
#define DESKTOP_ENUMERATE 0x0040L
#define DESKTOP_WRITEOBJECTS 0x0080L
#define DESKTOP_SWITCHDESKTOP 0x0100L
#define DF_ALLOWOTHERACCOUNTHOOK 0x0001L
#define WINSTA_ENUMDESKTOPS 0x0001L
#define WINSTA_READATTRIBUTES 0x0002L
#define WINSTA_ACCESSCLIPBOARD 0x0004L
#define WINSTA_CREATEDESKTOP 0x0008L
#define WINSTA_WRITEATTRIBUTES 0x0010L
#define WINSTA_ACCESSGLOBALATOMS 0x0020L
#define WINSTA_EXITWINDOWS 0x0040L
#define WINSTA_ENUMERATE 0x0100L
#define WINSTA_READSCREEN 0x0200L
#define WSF_VISIBLE 0x0001L
#define UOI_FLAGS 1
#define UOI_NAME 2
#define UOI_TYPE 3
#define GWL_WNDPROC (-4)
#define GWL_HINSTANCE (-6)
#define GWL_HWNDPARENT (-8)
#define GWL_STYLE (-16)
#define GWL_EXSTYLE (-20)
#define GWL_USERDATA (-21)
#define GWL_ID (-12)
#define GCL_MENUNAME (-8)
#define GCL_HBRBACKGROUND (-10)
#define GCL_HCURSOR (-12)
#define GCL_HICON (-14)
#define GCL_HMODULE (-16)
#define GCL_CBWNDEXTRA (-18)
#define GCL_CBCLSEXTRA (-20)
#define GCL_WNDPROC (-24)
#define GCL_STYLE (-26)
#define GCW_ATOM (-32)
#define GCL_HICONSM (-34)
#define WM_NULL 0x0000
#define WM_CREATE 0x0001
#define WM_DESTROY 0x0002
#define WM_MOVE 0x0003
#define WM_SIZE 0x0005
#define WM_ACTIVATE 0x0006
#define WA_INACTIVE 0
#define WA_ACTIVE 1
#define WA_CLICKACTIVE 2
#define WM_SETFOCUS 0x0007
#define WM_KILLFOCUS 0x0008
#define WM_ENABLE 0x000A
#define WM_SETREDRAW 0x000B
#define WM_SETTEXT 0x000C
#define WM_GETTEXT 0x000D
#define WM_GETTEXTLENGTH 0x000E
#define WM_PAINT 0x000F
#define WM_CLOSE 0x0010
#define WM_QUERYENDSESSION 0x0011
#define WM_QUIT 0x0012
#define WM_QUERYOPEN 0x0013
#define WM_ERASEBKGND 0x0014
#define WM_SYSCOLORCHANGE 0x0015
#define WM_ENDSESSION 0x0016
#define WM_SYSTEMERROR 0x0017
#define WM_SHOWWINDOW 0x0018
#define WM_CTLCOLOR 0x0019
#define WM_WININICHANGE 0x001A
#define WM_SETTINGCHANGE WM_WININICHANGE
#define WM_DEVMODECHANGE 0x001B
#define WM_ACTIVATEAPP 0x001C
#define WM_FONTCHANGE 0x001D
#define WM_TIMECHANGE 0x001E
#define WM_CANCELMODE 0x001F
#define WM_SETCURSOR 0x0020
#define WM_MOUSEACTIVATE 0x0021
#define WM_CHILDACTIVATE 0x0022
#define WM_QUEUESYNC 0x0023
#define WM_GETMINMAXINFO 0x0024
#define WM_PAINTICON 0x0026
#define WM_ICONERASEBKGND 0x0027
#define WM_NEXTDLGCTL 0x0028
#define WM_SPOOLERSTATUS 0x002A
#define WM_SETFONT 0x0030
#define WM_GETFONT 0x0031
#define WM_SETHOTKEY 0x0032
#define WM_GETHOTKEY 0x0033
#define WM_QUERYDRAGICON 0x0037
#define WM_GETOBJECT 0x003D
#define WM_COMPACTING 0x0041
#define WM_COMMNOTIFY 0x0044
#define WM_WINDOWPOSCHANGING 0x0046
#define WM_WINDOWPOSCHANGED 0x0047
#define WM_POWER 0x0048
#define PWR_OK 1
#define PWR_FAIL (-1)
#define PWR_SUSPENDREQUEST 1
#define PWR_SUSPENDRESUME 2
#define PWR_CRITICALRESUME 3
#define WM_COPYDATA 0x004A
#define WM_CANCELJOURNAL 0x004B
#define WM_NOTIFY 0x004E
#define WM_INPUTLANGCHANGEREQUEST 0x0050
#define WM_INPUTLANGCHANGE 0x0051
#define WM_TCARD 0x0052
#define WM_HELP 0x0053
#define WM_USERCHANGED 0x0054
#define WM_NOTIFYFORMAT 0x0055
#define NFR_ANSI 1
#define NFR_UNICODE 2
#define NF_QUERY 3
#define NF_REQUERY 4
#define WM_CONTEXTMENU 0x007B
#define WM_STYLECHANGING 0x007C
#define WM_STYLECHANGED 0x007D
#define WM_DISPLAYCHANGE 0x007E
#define WM_GETICON 0x007F
#define WM_SETICON 0x0080
#define WM_NCCREATE 0x0081
#define WM_NCDESTROY 0x0082
#define WM_NCCALCSIZE 0x0083
#define WM_NCHITTEST 0x0084
#define WM_NCPAINT 0x0085
#define WM_NCACTIVATE 0x0086
#define WM_GETDLGCODE 0x0087
#define WM_SYNCPAINT 0x0088
#define WM_NCMOUSEMOVE 0x00A0
#define WM_NCLBUTTONDOWN 0x00A1
#define WM_NCLBUTTONUP 0x00A2
#define WM_NCLBUTTONDBLCLK 0x00A3
#define WM_NCRBUTTONDOWN 0x00A4
#define WM_NCRBUTTONUP 0x00A5
#define WM_NCRBUTTONDBLCLK 0x00A6
#define WM_NCMBUTTONDOWN 0x00A7
#define WM_NCMBUTTONUP 0x00A8
#define WM_NCMBUTTONDBLCLK 0x00A9
#define WM_NCXBUTTONDOWN 0x00AB
#define WM_NCXBUTTONUP 0x00AC
#define WM_NCXBUTTONDBLCLK 0x00AD
#define WM_INPUT 0x00FF
#define WM_KEYFIRST 0x0100
#define WM_KEYDOWN 0x0100
#define WM_KEYUP 0x0101
#define WM_CHAR 0x0102
#define WM_DEADCHAR 0x0103
#define WM_SYSKEYDOWN 0x0104
#define WM_SYSKEYUP 0x0105
#define WM_SYSCHAR 0x0106
#define WM_SYSDEADCHAR 0x0107
#define WM_UNICHAR 0x0109
#define WM_KEYLAST 0x0109
#define UNICODE_NOCHAR 0xFFFF
#define WM_IME_STARTCOMPOSITION 0x010D
#define WM_IME_ENDCOMPOSITION 0x010E
#define WM_IME_COMPOSITION 0x010F
#define WM_IME_KEYLAST 0x010F
#define WM_INITDIALOG 0x0110
#define WM_SYSCOMMAND 0x0112
#define WM_TIMER 0x0113
#define WM_INITMENU 0x0116
#define WM_INITMENUPOPUP 0x0117
#define WM_SYSTIMER 0x0118U
#define WM_MENUSELECT 0x011F
#define WM_MENUCHAR 0x0120
#define WM_ENTERIDLE 0x0121
#define WM_MENURBUTTONUP 0x0122
#define WM_MENUDRAG 0x0123
#define WM_MENUGETOBJECT 0x0124
#define WM_UNINITMENUPOPUP 0x0125
#define WM_MENUCOMMAND 0x0126
#define WM_CHANGEUISTATE 0x0127
#define WM_UPDATEUISTATE 0x0128
#define WM_QUERYUISTATE 0x0129
#define UIS_SET 1
#define UIS_CLEAR 2
#define UIS_INITIALIZE 3
#define UISF_HIDEFOCUS 0x1
#define UISF_HIDEACCEL 0x2
#define UISF_ACTIVE 0x4
#define MN_GETHMENU 0x01E1
#define WM_MOUSEFIRST 0x0200
#define WM_MOUSEMOVE 0x0200
#define WM_LBUTTONDOWN 0x0201
#define WM_LBUTTONUP 0x0202
#define WM_LBUTTONDBLCLK 0x0203
#define WM_RBUTTONDOWN 0x0204
#define WM_RBUTTONUP 0x0205
#define WM_RBUTTONDBLCLK 0x0206
#define WM_MBUTTONDOWN 0x0207
#define WM_MBUTTONUP 0x0208
#define WM_MBUTTONDBLCLK 0x0209
#define WM_MOUSEWHEEL 0x020A
#define WM_XBUTTONDOWN 0x020B
#define WM_XBUTTONUP 0x020C
#define WM_XBUTTONDBLCLK 0x020D
#define WM_MOUSELAST 0x020D
#define WHEEL_DELTA 120
#define WHEEL_PAGESCROLL (0xFFFFFFFF)
#define MENULOOP_WINDOW 0
#define MENULOOP_POPUP 1
#define WM_ENTERMENULOOP 0x0211
#define WM_EXITMENULOOP 0x0212
#define WM_NEXTMENU 0x0213
#define WM_SIZING 0x0214
#define WM_CAPTURECHANGED 0x0215
#define WM_MOVING 0x0216
#define WM_POWERBROADCAST 0x0218
#define WM_DEVICECHANGE 0x0219
#define WM_MDICREATE 0x0220
#define WM_MDIDESTROY 0x0221
#define WM_MDIACTIVATE 0x0222
#define WM_MDIRESTORE 0x0223
#define WM_MDINEXT 0x0224
#define WM_MDIMAXIMIZE 0x0225
#define WM_MDITILE 0x0226
#define WM_MDICASCADE 0x0227
#define WM_MDIICONARRANGE 0x0228
#define WM_MDIGETACTIVE 0x0229
#define WM_MDISETMENU 0x0230
#define WM_ENTERSIZEMOVE 0x0231
#define WM_EXITSIZEMOVE 0x0232
#define WM_DROPFILES 0x0233
#define WM_MDIREFRESHMENU 0x0234
#define WM_IME_SETCONTEXT 0x0281
#define WM_IME_NOTIFY 0x0282
#define WM_IME_CONTROL 0x0283
#define WM_IME_COMPOSITIONFULL 0x0284
#define WM_IME_SELECT 0x0285
#define WM_IME_CHAR 0x0286
#define WM_IME_REQUEST 0x0288
#define WM_IME_KEYDOWN 0x0290
#define WM_IME_KEYUP 0x0291
#define WM_MOUSEHOVER 0x02A1
#define WM_MOUSELEAVE 0x02A3
#define WM_NCMOUSEHOVER 0x02A0
#define WM_NCMOUSELEAVE 0x02A2
#define WM_WTSSESSION_CHANGE 0x02B1
#define WM_TABLET_FIRST 0x02c0
#define WM_TABLET_LAST 0x02df
#define WM_CUT 0x0300
#define WM_COPY 0x0301
#define WM_PASTE 0x0302
#define WM_CLEAR 0x0303
#define WM_UNDO 0x0304
#define WM_RENDERFORMAT 0x0305
#define WM_RENDERALLFORMATS 0x0306
#define WM_DESTROYCLIPBOARD 0x0307
#define WM_DRAWCLIPBOARD 0x0308
#define WM_PAINTCLIPBOARD 0x0309
#define WM_VSCROLLCLIPBOARD 0x030A
#define WM_SIZECLIPBOARD 0x030B
#define WM_ASKCBFORMATNAME 0x030C
#define WM_CHANGECBCHAIN 0x030D
#define WM_HSCROLLCLIPBOARD 0x030E
#define WM_QUERYNEWPALETTE 0x030F
#define WM_PALETTEISCHANGING 0x0310
#define WM_PALETTECHANGED 0x0311
#define WM_HOTKEY 0x0312
#define WM_PRINT 0x0317
#define WM_PRINTCLIENT 0x0318
#define WM_APPCOMMAND 0x0319
#define WM_THEMECHANGED 0x031A
#define WM_HANDHELDFIRST 0x0358
#define WM_HANDHELDLAST 0x035F
#define WM_AFXFIRST 0x0360
#define WM_AFXLAST 0x037F
#define WM_PENWINFIRST 0x0380
#define WM_PENWINLAST 0x038F
#define WM_APP 0x8000
#define WM_VOAPP WM_APP + 0x1000
#define WMSZ_LEFT 1
#define WMSZ_RIGHT 2
#define WMSZ_TOP 3
#define WMSZ_TOPLEFT 4
#define WMSZ_TOPRIGHT 5
#define WMSZ_BOTTOM 6
#define WMSZ_BOTTOMLEFT 7
#define WMSZ_BOTTOMRIGHT 8
#define ST_BEGINSWP 0
#define ST_ENDSWP 1
#define HTERROR (-2)
#define HTTRANSPARENT (-1)
#define HTNOWHERE 0
#define HTCLIENT 1
#define HTCAPTION 2
#define HTSYSMENU 3
#define HTGROWBOX 4
#define HTSIZE HTGROWBOX
#define HTMENU 5
#define HTHSCROLL 6
#define HTVSCROLL 7
#define HTMINBUTTON 8
#define HTMAXBUTTON 9
#define HTLEFT 10
#define HTRIGHT 11
#define HTTOP 12
#define HTTOPLEFT 13
#define HTTOPRIGHT 14
#define HTBOTTOM 15
#define HTBOTTOMLEFT 16
#define HTBOTTOMRIGHT 17
#define HTBORDER 18
#define HTREDUCE HTMINBUTTON
#define HTZOOM HTMAXBUTTON
#define HTSIZEFIRST HTLEFT
#define HTSIZELAST HTBOTTOMRIGHT
#define HTOBJECT 19
#define HTCLOSE 20
#define HTHELP 21
#define SMTO_NORMAL 0x0000
#define SMTO_BLOCK 0x0001
#define SMTO_ABORTIFHUNG 0x0002
#define SMTO_NOTIMEOUTIFNOTHUNG 0x0008
#define MA_ACTIVATE 1
#define MA_ACTIVATEANDEAT 2
#define MA_NOACTIVATE 3
#define MA_NOACTIVATEANDEAT 4
#define ICON_SMALL 0
#define ICON_BIG 1
#define SIZE_RESTORED 0
#define SIZE_MINIMIZED 1
#define SIZE_MAXIMIZED 2
#define SIZE_MAXSHOW 3
#define SIZE_MAXHIDE 4
#define SIZENORMAL SIZE_RESTORED
#define SIZEICONIC SIZE_MINIMIZED
#define SIZEFULLSCREEN SIZE_MAXIMIZED
#define SIZEZOOMSHOW SIZE_MAXSHOW
#define SIZEZOOMHIDE SIZE_MAXHIDE
#define WVR_ALIGNTOP 0x0010
#define WVR_ALIGNLEFT 0x0020
#define WVR_ALIGNBOTTOM 0x0040
#define WVR_ALIGNRIGHT 0x0080
#define WVR_HREDRAW 0x0100
#define WVR_VREDRAW 0x0200
#define WVR_REDRAW 0x0300
#define WVR_VALIDRECTS 0x0400
#define MK_LBUTTON 0x0001
#define MK_RBUTTON 0x0002
#define MK_SHIFT 0x0004
#define MK_CONTROL 0x0008
#define MK_MBUTTON 0x0010
#define MK_XBUTTON1 0x0020
#define MK_XBUTTON2 0x0040
#define WS_OVERLAPPED 0x00000000L
#define WS_POPUP 0x80000000
#define WS_CHILD 0x40000000L
#define WS_MINIMIZE 0x20000000L
#define WS_VISIBLE 0x10000000L
#define WS_DISABLED 0x08000000L
#define WS_CLIPSIBLINGS 0x04000000L
#define WS_CLIPCHILDREN 0x02000000L
#define WS_MAXIMIZE 0x01000000L
#define WS_CAPTION 0x00C00000L
#define WS_BORDER 0x00800000L
#define WS_DLGFRAME 0x00400000L
#define WS_VSCROLL 0x00200000L
#define WS_HSCROLL 0x00100000L
#define WS_SYSMENU 0x00080000L
#define WS_THICKFRAME 0x00040000L
#define WS_GROUP 0x00020000L
#define WS_TABSTOP 0x00010000L
#define WS_MINIMIZEBOX 0x00020000L
#define WS_MAXIMIZEBOX 0x00010000L
#define WS_TILED WS_OVERLAPPED
#define WS_ICONIC WS_MINIMIZE
#define WS_SIZEBOX WS_THICKFRAME
#define WS_OVERLAPPEDWINDOW 0x00CF0000L
#define WS_TILEDWINDOW WS_OVERLAPPEDWINDOW
#define WS_POPUPWINDOW 0X80880000
#define WS_CHILDWINDOW (WS_CHILD)
#define WS_EX_DLGMODALFRAME 0x00000001L
#define WS_EX_NOPARENTNOTIFY 0x00000004L
#define WS_EX_TOPMOST 0x00000008L
#define WS_EX_ACCEPTFILES 0x00000010L
#define WS_EX_TRANSPARENT 0x00000020L
#define WS_EX_MDICHILD 0x00000040L
#define WS_EX_TOOLWINDOW 0x00000080L
#define WS_EX_WINDOWEDGE 0x00000100L
#define WS_EX_CLIENTEDGE 0x00000200L
#define WS_EX_CONTEXTHELP 0x00000400L
#define WS_EX_RIGHT 0x00001000L
#define WS_EX_LEFT 0x00000000L
#define WS_EX_RTLREADING 0x00002000L
#define WS_EX_LTRREADING 0x00000000L
#define WS_EX_LEFTSCROLLBAR 0x00004000L
#define WS_EX_RIGHTSCROLLBAR 0x00000000L
#define WS_EX_CONTROLPARENT 0x00010000L
#define WS_EX_STATICEDGE 0x00020000L
#define WS_EX_APPWINDOW 0x00040000L
#define WS_EX_OVERLAPPEDWINDOW 0x00000300L
#define WS_EX_PALETTEWINDOW 0x00000188L
#define WS_EX_LAYERED 0x00080000
#define WS_EX_NOINHERITLAYOUT 0x00100000L
#define WS_EX_LAYOUTRTL 0x00400000L
#define CS_VREDRAW 0x0001
#define CS_HREDRAW 0x0002
#define CS_KEYCVTWINDOW 0x0004
#define CS_DBLCLKS 0x0008
#define CS_OWNDC 0x0020
#define CS_CLASSDC 0x0040
#define CS_PARENTDC 0x0080
#define CS_NOKEYCVT 0x0100
#define CS_NOCLOSE 0x0200
#define CS_SAVEBITS 0x0800
#define CS_BYTEALIGNCLIENT 0x1000
#define CS_BYTEALIGNWINDOW 0x2000
#define CS_GLOBALCLASS 0x4000
#define CS_IME 0x00010000
#define CS_DROPSHADOW 0x00020000
#define PRF_CHECKVISIBLE 0x00000001L
#define PRF_NONCLIENT 0x00000002L
#define PRF_CLIENT 0x00000004L
#define PRF_ERASEBKGND 0x00000008L
#define PRF_CHILDREN 0x00000010L
#define PRF_OWNED 0x00000020L
#define BDR_RAISEDOUTER 0x0001
#define BDR_SUNKENOUTER 0x0002
#define BDR_RAISEDINNER 0x0004
#define BDR_SUNKENINNER 0x0008
#define BDR_OUTER 0x0003
#define BDR_INNER 0x000c
#define BDR_RAISED 0x0005
#define BDR_SUNKEN 0x000a
#define EDGE_RAISED 0x0005
#define EDGE_SUNKEN 0x000A
#define EDGE_ETCHED 0x0006
#define EDGE_BUMP 0x0009
#define BF_LEFT 0x0001
#define BF_TOP 0x0002
#define BF_RIGHT 0x0004
#define BF_BOTTOM 0x0008
#define BF_TOPLEFT 0x0003
#define BF_TOPRIGHT 0x0006
#define BF_BOTTOMLEFT 0x0009
#define BF_BOTTOMRIGHT 0x000C
#define BF_RECT 0x000F
#define BF_DIAGONAL 0x0010
#define BF_DIAGONAL_ENDTOPRIGHT 0x0016
#define BF_DIAGONAL_ENDTOPLEFT 0x0013
#define BF_DIAGONAL_ENDBOTTOMLEFT 0x0019
#define BF_DIAGONAL_ENDBOTTOMRIGHT 0x001C
#define BF_MIDDLE 0x0800
#define BF_SOFT 0x1000
#define BF_ADJUST 0x2000
#define BF_FLAT 0x4000
#define BF_MONO 0x8000
#define DFC_CAPTION 1
#define DFC_MENU 2
#define DFC_SCROLL 3
#define DFC_BUTTON 4
#define DFC_POPUPMENU 5
#define DFCS_CAPTIONCLOSE 0x0000
#define DFCS_CAPTIONMIN 0x0001
#define DFCS_CAPTIONMAX 0x0002
#define DFCS_CAPTIONRESTORE 0x0003
#define DFCS_CAPTIONHELP 0x0004
#define DFCS_MENUARROW 0x0000
#define DFCS_MENUCHECK 0x0001
#define DFCS_MENUBULLET 0x0002
#define DFCS_MENUARROWRIGHT 0x0004
#define DFCS_SCROLLUP 0x0000
#define DFCS_SCROLLDOWN 0x0001
#define DFCS_SCROLLLEFT 0x0002
#define DFCS_SCROLLRIGHT 0x0003
#define DFCS_SCROLLCOMBOBOX 0x0005
#define DFCS_SCROLLSIZEGRIP 0x0008
#define DFCS_SCROLLSIZEGRIPRIGHT 0x0010
#define DFCS_BUTTONCHECK 0x0000
#define DFCS_BUTTONRADIOIMAGE 0x0001
#define DFCS_BUTTONRADIOMASK 0x0002
#define DFCS_BUTTONRADIO 0x0004
#define DFCS_BUTTON3STATE 0x0008
#define DFCS_BUTTONPUSH 0x0010
#define DFCS_INACTIVE 0x0100
#define DFCS_PUSHED 0x0200
#define DFCS_CHECKED 0x0400
#define DFCS_TRANSPARENT 0x0800
#define DFCS_HOT 0x1000
#define DFCS_ADJUSTRECT 0x2000
#define DFCS_FLAT 0x4000
#define DFCS_MONO 0x8000
#define DC_ACTIVE 0x0001
#define DC_SMALLCAP 0x0002
#define DC_ICON 0x0004
#define DC_TEXT 0x0008
#define DC_INBUTTON 0x0010
#define DC_GRADIENT 0x0020
#define DC_BUTTONS 0x1000
#define IDANI_OPEN 1
#define IDANI_CLOSE 2
#define IDANI_CAPTION 3
#define CF_TEXT 1
#define CF_BITMAP 2
#define CF_METAFILEPICT 3
#define CF_SYLK 4
#define CF_DIF 5
#define CF_TIFF 6
#define CF_OEMTEXT 7
#define CF_DIB 8
#define CF_PALETTE 9
#define CF_PENDATA 10
#define CF_RIFF 11
#define CF_WAVE 12
#define CF_UNICODETEXT 13
#define CF_ENHMETAFILE 14
#define CF_HDROP 15
#define CF_LOCALE 16
#define CF_DIBV5 17
#define CF_MAX 17
#define CF_OWNERDISPLAY 0x0080
#define CF_DSPTEXT 0x0081
#define CF_DSPBITMAP 0x0082
#define CF_DSPMETAFILEPICT 0x0083
#define CF_DSPENHMETAFILE 0x008E
#define CF_PRIVATEFIRST 0x0200
#define CF_PRIVATELAST 0x02FF
#define CF_GDIOBJFIRST 0x0300
#define CF_GDIOBJLAST 0x03FF
#define FVIRTKEY TRUE
#define FNOINVERT 0x02
#define FSHIFT 0x04
#define FCONTROL 0x08
#define FALT 0x10
#define WPF_SETMINPOSITION 0x0001
#define WPF_RESTORETOMAXIMIZED 0x0002
#define ODT_MENU 1
#define ODT_LISTBOX 2
#define ODT_COMBOBOX 3
#define ODT_BUTTON 4
#define ODT_STATIC 5
#define ODA_DRAWENTIRE 0x0001
#define ODA_SELECT 0x0002
#define ODA_FOCUS 0x0004
#define ODS_SELECTED 0x0001
#define ODS_GRAYED 0x0002
#define ODS_DISABLED 0x0004
#define ODS_CHECKED 0x0008
#define ODS_FOCUS 0x0010
#define ODS_DEFAULT 0x0020
#define ODS_COMBOBOXEDIT 0x1000
#define ODS_HOTLIGHT 0x0040
#define ODS_INACTIVE 0x0080
#define ODS_NOACCEL 0x0100
#define ODS_NOFOCUSRECT 0x0200
#define PM_NOREMOVE 0x0000
#define PM_REMOVE 0x0001
#define PM_NOYIELD 0x0002
#define MOD_ALT 0x0001
#define MOD_CONTROL 0x0002
#define MOD_SHIFT 0x0004
#define MOD_WIN 0x0008
#define IDHOT_SNAPWINDOW (-1)
#define IDHOT_SNAPDESKTOP (-2)
#define EW_RESTARTWINDOWS 0x0042L
#define EW_REBOOTSYSTEM 0x0043L
#define EW_EXITANDEXECAPP 0x0044L
#define EWX_LOGOFF 0
#define EWX_SHUTDOWN 1
#define EWX_REBOOT 2
#define EWX_FORCE 4
#define EWX_POWEROFF 8
#define EWX_FORCEIFHUNG 0x00000010
#define BSM_ALLCOMPONENTS 0x00000000
#define BSM_VXDS 0x00000001
#define BSM_NETDRIVER 0x00000002
#define BSM_INSTALLABLEDRIVERS 0x00000004
#define BSM_APPLICATIONS 0x00000008
#define BSM_ALLDESKTOPS 0x00000010
#define BSF_QUERY 0x00000001
#define BSF_IGNORECURRENTTASK 0x00000002
#define BSF_FLUSHDISK 0x00000004
#define BSF_NOHANG 0x00000008
#define BSF_POSTMESSAGE 0x00000010
#define BSF_FORCEIFHUNG 0x00000020
#define BSF_NOTIMEOUTIFNOTHUNG 0x00000040
#define BSF_ALLOWSFW 0x00000080
#define BSF_SENDNOTIFYMESSAGE 0x00000100
#define BSF_RETURNHDESK 0x00000200
#define BSF_LUID 0x00000400
#define DBWF_LPARAMPOINTER 0x8000
#define BROADCAST_QUERY_DENY 0x424D5144
#define HWND_BROADCAST PTR(_CAST, 0xffff)
#define CW_USEDEFAULT INT(_CAST,0x80000000)
#define HWND_DESKTOP PTR(_CAST, 0)
#define SWP_NOSIZE 0x0001
#define SWP_NOMOVE 0x0002
#define SWP_NOZORDER 0x0004
#define SWP_NOREDRAW 0x0008
#define SWP_NOACTIVATE 0x0010
#define SWP_FRAMECHANGED 0x0020
#define SWP_SHOWWINDOW 0x0040
#define SWP_HIDEWINDOW 0x0080
#define SWP_NOCOPYBITS 0x0100
#define SWP_NOOWNERZORDER 0x0200
#define SWP_NOSENDCHANGING 0x0400
#define SWP_DRAWFRAME SWP_FRAMECHANGED
#define SWP_NOREPOSITION SWP_NOOWNERZORDER
#define SWP_DEFERERASE 0x2000
#define SWP_ASYNCWINDOWPOS 0x4000
#define HWND_TOP PTR(_CAST, 0)
#define HWND_BOTTOM PTR(_CAST, 1)
#define HWND_TOPMOST PTR(_CAST, 0xFFFFFFFF)
#define HWND_NOTOPMOST PTR(_CAST, 0xFFFFFFFE)
#define DLGWINDOWEXTRA 30
#define KEYEVENTF_EXTENDEDKEY 0x0001
#define KEYEVENTF_KEYUP 0x0002
#define MOUSEEVENTF_MOVE 0x0001
#define MOUSEEVENTF_LEFTDOWN 0x0002
#define MOUSEEVENTF_LEFTUP 0x0004
#define MOUSEEVENTF_RIGHTDOWN 0x0008
#define MOUSEEVENTF_RIGHTUP 0x0010
#define MOUSEEVENTF_MIDDLEDOWN 0x0020
#define MOUSEEVENTF_MIDDLEUP 0x0040
#define MOUSEEVENTF_XDOWN 0x0080 
#define MOUSEEVENTF_XUP 0x0100 
#define MOUSEEVENTF_WHEEL 0x0800 
#define MOUSEEVENTF_VIRTUALDESK 0x4000 
#define MOUSEEVENTF_ABSOLUTE 0x8000
#define QS_KEY 0x0001
#define QS_MOUSEMOVE 0x0002
#define QS_MOUSEBUTTON 0x0004
#define QS_POSTMESSAGE 0x0008
#define QS_TIMER 0x0010
#define QS_PAINT 0x0020
#define QS_SENDMESSAGE 0x0040
#define QS_HOTKEY 0x0080
#define QS_ALLPOSTMESSAGE 0x0100
#define QS_RAWINPUT 0x0400
#define QS_MOUSE 0x0006
#define QS_INPUT 0x0007
#define QS_ALLEVENTS 0x00BF
#define QS_ALLINPUT 0x00FF
#define USER_TIMER_MAXIMUM 0x7FFFFFFF
#define USER_TIMER_MINIMUM 0x0000000A
#define SM_CXSCREEN 0
#define SM_CYSCREEN 1
#define SM_CXVSCROLL 2
#define SM_CYHSCROLL 3
#define SM_CYCAPTION 4
#define SM_CXBORDER 5
#define SM_CYBORDER 6
#define SM_CXDLGFRAME 7
#define SM_CYDLGFRAME 8
#define SM_CYVTHUMB 9
#define SM_CXHTHUMB 10
#define SM_CXICON 11
#define SM_CYICON 12
#define SM_CXCURSOR 13
#define SM_CYCURSOR 14
#define SM_CYMENU 15
#define SM_CXFULLSCREEN 16
#define SM_CYFULLSCREEN 17
#define SM_CYKANJIWINDOW 18
#define SM_MOUSEPRESENT 19
#define SM_CYVSCROLL 20
#define SM_CXHSCROLL 21
#define SM_DEBUG 22
#define SM_SWAPBUTTON 23
#define SM_RESERVED1 24
#define SM_RESERVED2 25
#define SM_RESERVED3 26
#define SM_RESERVED4 27
#define SM_CXMIN 28
#define SM_CYMIN 29
#define SM_CXSIZE 30
#define SM_CYSIZE 31
#define SM_CXFRAME 32
#define SM_CYFRAME 33
#define SM_CXMINTRACK 34
#define SM_CYMINTRACK 35
#define SM_CXDOUBLECLK 36
#define SM_CYDOUBLECLK 37
#define SM_CXICONSPACING 38
#define SM_CYICONSPACING 39
#define SM_MENUDROPALIGNMENT 40
#define SM_PENWINDOWS 41
#define SM_DBCSENABLED 42
#define SM_CMOUSEBUTTONS 43
#define SM_CXFIXEDFRAME SM_CXDLGFRAME
#define SM_CYFIXEDFRAME SM_CYDLGFRAME
#define SM_CXSIZEFRAME SM_CXFRAME
#define SM_CYSIZEFRAME SM_CYFRAME
#define SM_SECURE 44
#define SM_CXEDGE 45
#define SM_CYEDGE 46
#define SM_CXMINSPACING 47
#define SM_CYMINSPACING 48
#define SM_CXSMICON 49
#define SM_CYSMICON 50
#define SM_CYSMCAPTION 51
#define SM_CXSMSIZE 52
#define SM_CYSMSIZE 53
#define SM_CXMENUSIZE 54
#define SM_CYMENUSIZE 55
#define SM_ARRANGE 56
#define SM_CXMINIMIZED 57
#define SM_CYMINIMIZED 58
#define SM_CXMAXTRACK 59
#define SM_CYMAXTRACK 60
#define SM_CXMAXIMIZED 61
#define SM_CYMAXIMIZED 62
#define SM_NETWORK 63
#define SM_CLEANBOOT 67
#define SM_CXDRAG 68
#define SM_CYDRAG 69
#define SM_SHOWSOUNDS 70
#define SM_CXMENUCHECK 71
#define SM_CYMENUCHECK 72
#define SM_SLOWMACHINE 73
#define SM_MIDEASTENABLED 74
#define SM_MOUSEWHEELPRESENT 75
#define SM_XVIRTUALSCREEN 76
#define SM_YVIRTUALSCREEN 77
#define SM_CXVIRTUALSCREEN 78
#define SM_CYVIRTUALSCREEN 79
#define SM_CMONITORS 80
#define SM_SAMEDISPLAYFORMAT 81
#define SM_IMMENABLED 82
#define SM_CXFOCUSBORDER 83
#define SM_CYFOCUSBORDER 84
#define SM_TABLETPC 86
#define SM_MEDIACENTER 87
#define SM_STARTER 88
#define SM_SERVERR2 89
#define SM_REMOTESESSION 0x1000
#define SM_SHUTTINGDOWN 0x2000
#define SM_REMOTECONTROL 0x2001
#define SM_CARETBLINKINGENABLED 0x2002
#define MNC_IGNORE 0
#define MNC_CLOSE 1
#define MNC_EXECUTE 2
#define MNC_SELECT 3
#define MIIM_STATE 0x00000001
#define MIIM_ID 0x00000002
#define MIIM_SUBMENU 0x00000004
#define MIIM_CHECKMARKS 0x00000008
#define MIIM_TYPE 0x00000010
#define MIIM_DATA 0x00000020
#define GMDI_USEDISABLED 0x0001L
#define GMDI_GOINTOPOPUPS 0x0002L
#define TPM_LEFTBUTTON 0x0000L
#define TPM_RIGHTBUTTON 0x0002L
#define TPM_LEFTALIGN 0x0000L
#define TPM_CENTERALIGN 0x0004L
#define TPM_RIGHTALIGN 0x0008L
#define TPM_TOPALIGN 0x0000L
#define TPM_VCENTERALIGN 0x0010L
#define TPM_BOTTOMALIGN 0x0020L
#define TPM_HORIZONTAL 0x0000L
#define TPM_VERTICAL 0x0040L
#define TPM_NONOTIFY 0x0080L
#define TPM_RETURNCMD 0x0100L
#define DOF_EXECUTABLE 0x8001
#define DOF_DOCUMENT 0x8002
#define DOF_DIRECTORY 0x8003
#define DOF_MULTIPLE 0x8004
#define DOF_PROGMAN 0x0001
#define DOF_SHELLDATA 0x0002
#define DO_DROPFILE 0x454C4946L
#define DO_PRINTFILE 0x544E5250L
#define DT_TOP 0x00000000
#define DT_LEFT 0x00000000
#define DT_CENTER 0x00000001
#define DT_RIGHT 0x00000002
#define DT_VCENTER 0x00000004
#define DT_BOTTOM 0x00000008
#define DT_WORDBREAK 0x00000010
#define DT_SINGLELINE 0x00000020
#define DT_EXPANDTABS 0x00000040
#define DT_TABSTOP 0x00000080
#define DT_NOCLIP 0x00000100
#define DT_EXTERNALLEADING 0x00000200
#define DT_CALCRECT 0x00000400
#define DT_NOPREFIX 0x00000800
#define DT_INTERNAL 0x00001000
#define DT_EDITCONTROL 0x00002000
#define DT_PATH_ELLIPSIS 0x00004000
#define DT_END_ELLIPSIS 0x00008000
#define DT_MODIFYSTRING 0x00010000
#define DT_RTLREADING 0x00020000
#define DT_WORD_ELLIPSIS 0x00040000
#define DST_COMPLEX 0x0000
#define DST_TEXT 0x0001
#define DST_PREFIXTEXT 0x0002
#define DST_ICON 0x0003
#define DST_BITMAP 0x0004
#define DSS_NORMAL 0x0000
#define DSS_UNION 0x0010
#define DSS_DISABLED 0x0020
#define DSS_MONO 0x0080
#define DSS_RIGHT 0x8000
#define DCX_WINDOW 0x00000001L
#define DCX_CACHE 0x00000002L
#define DCX_NORESETATTRS 0x00000004L
#define DCX_CLIPCHILDREN 0x00000008L
#define DCX_CLIPSIBLINGS 0x00000010L
#define DCX_PARENTCLIP 0x00000020L
#define DCX_EXCLUDERGN 0x00000040L
#define DCX_INTERSECTRGN 0x00000080L
#define DCX_EXCLUDEUPDATE 0x00000100L
#define DCX_INTERSECTUPDATE 0x00000200L
#define DCX_LOCKWINDOWUPDATE 0x00000400L
#define DCX_VALIDATE 0x00200000L
#define RDW_INVALIDATE 0x0001
#define RDW_INTERNALPAINT 0x0002
#define RDW_ERASE 0x0004
#define RDW_VALIDATE 0x0008
#define RDW_NOINTERNALPAINT 0x0010
#define RDW_NOERASE 0x0020
#define RDW_NOCHILDREN 0x0040
#define RDW_ALLCHILDREN 0x0080
#define RDW_UPDATENOW 0x0100
#define RDW_ERASENOW 0x0200
#define RDW_FRAME 0x0400
#define RDW_NOFRAME 0x0800
#define SW_SCROLLCHILDREN 0x0001
#define SW_INVALIDATE 0x0002
#define SW_ERASE 0x0004
#define ESB_ENABLE_BOTH 0x0000
#define ESB_DISABLE_BOTH 0x0003
#define ESB_DISABLE_LEFT 0x0001
#define ESB_DISABLE_RIGHT 0x0002
#define ESB_DISABLE_UP 0x0001
#define ESB_DISABLE_DOWN 0x0002
#define ESB_DISABLE_LTUP ESB_DISABLE_LEFT
#define ESB_DISABLE_RTDN ESB_DISABLE_RIGHT
#define HELPINFO_WINDOW 0x0001
#define HELPINFO_MENUITEM 0x0002
#define MB_OK 0x00000000U
#define MB_OKCANCEL 0x00000001U
#define MB_ABORTRETRYIGNORE 0x00000002U
#define MB_YESNOCANCEL 0x00000003U
#define MB_YESNO 0x00000004U
#define MB_RETRYCANCEL 0x00000005U
#define MB_CANCELTRYCONTINUE 0x00000006U
#define MB_ICONHAND 0x00000010U
#define MB_ICONQUESTION 0x00000020U
#define MB_ICONEXCLAMATION 0x00000030U
#define MB_ICONASTERISK 0x00000040U
#define MB_USERICON 0x00000080U
#define MB_ICONWARNING MB_ICONEXCLAMATION
#define MB_ICONERROR MB_ICONHAND
#define MB_ICONINFORMATION MB_ICONASTERISK
#define MB_ICONSTOP MB_ICONHAND
#define MB_DEFBUTTON1 0x00000000U
#define MB_DEFBUTTON2 0x00000100U
#define MB_DEFBUTTON3 0x00000200U
#define MB_DEFBUTTON4 0x00000300U
#define MB_APPLMODAL 0x00000000U
#define MB_SYSTEMMODAL 0x00001000U
#define MB_TASKMODAL 0x00002000U
#define MB_HELP 0x00004000U
#define MB_NOFOCUS 0x00008000U
#define MB_SETFOREGROUND 0x00010000U
#define MB_DEFAULT_DESKTOP_ONLY 0x00020000U
#define MB_TOPMOST 0x00040000U
#define MB_RIGHT 0x00080000U
#define MB_RTLREADING 0x00100000U
#define MB_SERVICE_NOTIFICATION 0x00040000U
#define MB_TYPEMASK 0x0000000FU
#define MB_ICONMASK 0x000000F0U
#define MB_DEFMASK 0x00000F00U
#define MB_MODEMASK 0x00003000U
#define MB_MISCMASK 0x0000C000U
#define CWP_ALL 0x0000
#define CWP_SKIPINVISIBLE 0x0001
#define CWP_SKIPDISABLED 0x0002
#define CWP_SKIPTRANSPARENT 0x0004
#define CTLCOLOR_MSGBOX 0
#define CTLCOLOR_EDIT 1
#define CTLCOLOR_LISTBOX 2
#define CTLCOLOR_BTN 3
#define CTLCOLOR_DLG 4
#define CTLCOLOR_SCROLLBAR 5
#define CTLCOLOR_STATIC 6
#define CTLCOLOR_MAX 7
#define COLOR_SCROLLBAR 0
#define COLOR_BACKGROUND 1
#define COLOR_ACTIVECAPTION 2
#define COLOR_INACTIVECAPTION 3
#define COLOR_MENU 4
#define COLOR_WINDOW 5
#define COLOR_WINDOWFRAME 6
#define COLOR_MENUTEXT 7
#define COLOR_WINDOWTEXT 8
#define COLOR_CAPTIONTEXT 9
#define COLOR_ACTIVEBORDER 10
#define COLOR_INACTIVEBORDER 11
#define COLOR_APPWORKSPACE 12
#define COLOR_HIGHLIGHT 13
#define COLOR_HIGHLIGHTTEXT 14
#define COLOR_BTNFACE 15
#define COLOR_BTNSHADOW 16
#define COLOR_GRAYTEXT 17
#define COLOR_BTNTEXT 18
#define COLOR_INACTIVECAPTIONTEXT 19
#define COLOR_BTNHIGHLIGHT 20
#define COLOR_3DDKSHADOW 21
#define COLOR_3DLIGHT 22
#define COLOR_INFOTEXT 23
#define COLOR_INFOBK 24
#define COLOR_HOTLIGHT 26
#define COLOR_GRADIENTACTIVECAPTION 27
#define COLOR_GRADIENTINACTIVECAPTION 28
#define COLOR_MENUHILIGHT 29
#define COLOR_MENUBAR 30
#define COLOR_DESKTOP COLOR_BACKGROUND
#define COLOR_3DFACE COLOR_BTNFACE
#define COLOR_3DSHADOW COLOR_BTNSHADOW
#define COLOR_3DHIGHLIGHT COLOR_BTNHIGHLIGHT
#define COLOR_3DHILIGHT COLOR_BTNHIGHLIGHT
#define COLOR_BTNHILIGHT COLOR_BTNHIGHLIGHT
#define GW_HWNDFIRST 0
#define GW_HWNDLAST 1
#define GW_HWNDNEXT 2
#define GW_HWNDPREV 3
#define GW_OWNER 4
#define GW_CHILD 5
#define GW_ENABLEDPOPUP 6
#define GW_MAX 6
#define MF_INSERT 0x00000000L
#define MF_CHANGE 0x00000080L
#define MF_APPEND 0x00000100L
#define MF_DELETE 0x00000200L
#define MF_REMOVE 0x00001000L
#define MF_BYCOMMAND 0x00000000L
#define MF_BYPOSITION 0x00000400L
#define MF_SEPARATOR 0x00000800L
#define MF_ENABLED 0x00000000L
#define MF_GRAYED 0x00000001L
#define MF_DISABLED 0x00000002L
#define MF_UNCHECKED 0x00000000L
#define MF_CHECKED 0x00000008L
#define MF_USECHECKBITMAPS 0x00000200L
#define MF_STRING 0x00000000L
#define MF_BITMAP 0x00000004L
#define MF_OWNERDRAW 0x00000100L
#define MF_POPUP 0x00000010L
#define MF_MENUBARBREAK 0x00000020L
#define MF_MENUBREAK 0x00000040L
#define MF_UNHILITE 0x00000000L
#define MF_HILITE 0x00000080L
#define MF_DEFAULT 0x00001000L
#define MF_SYSMENU 0x00002000L
#define MF_HELP 0x00004000L
#define MF_RIGHTJUSTIFY 0x00004000L
#define MF_MOUSESELECT 0x00008000L
#define MF_END 0x00000080L
#define MFT_STRING MF_STRING
#define MFT_BITMAP MF_BITMAP
#define MFT_MENUBARBREAK MF_MENUBARBREAK
#define MFT_MENUBREAK MF_MENUBREAK
#define MFT_OWNERDRAW MF_OWNERDRAW
#define MFT_RADIOCHECK 0x00000200L
#define MFT_SEPARATOR MF_SEPARATOR
#define MFT_RIGHTORDER 0x00002000L
#define MFT_RIGHTJUSTIFY MF_RIGHTJUSTIFY
#define MFS_GRAYED 0x00000003L
#define MFS_DISABLED MFS_GRAYED
#define MFS_CHECKED MF_CHECKED
#define MFS_HILITE MF_HILITE
#define MFS_ENABLED MF_ENABLED
#define MFS_UNCHECKED MF_UNCHECKED
#define MFS_UNHILITE MF_UNHILITE
#define MFS_DEFAULT MF_DEFAULT
#define SC_MOVE 0xF010
#define SC_MINIMIZE 0xF020
#define SC_MAXIMIZE 0xF030
#define SC_NEXTWINDOW 0xF040
#define SC_PREVWINDOW 0xF050
#define SC_CLOSE 0xF060
#define SC_VSCROLL 0xF070
#define SC_HSCROLL 0xF080
#define SC_MOUSEMENU 0xF090
#define SC_KEYMENU 0xF100
#define SC_ARRANGE 0xF110
#define SC_RESTORE 0xF120
#define SC_TASKLIST 0xF130
#define SC_SCREENSAVE 0xF140
#define SC_HOTKEY 0xF150
#define SC_DEFAULT 0xF160
#define SC_MONITORPOWER 0xF170
#define SC_CONTEXTHELP 0xF180
#define SC_SEPARATOR 0xF00F
#define SC_ICON SC_MINIMIZE
#define SC_ZOOM SC_MAXIMIZE
#define IDC_ARROW PTR(_CAST, 32512)
#define IDC_IBEAM PTR(_CAST, 32513)
#define IDC_WAIT PTR(_CAST, 32514)
#define IDC_CROSS PTR(_CAST, 32515)
#define IDC_UPARROW PTR(_CAST, 32516)
#define IDC_SIZE PTR(_CAST, 32640)
#define IDC_ICON PTR(_CAST, 32641)
#define IDC_SIZENWSE PTR(_CAST, 32642)
#define IDC_SIZENESW PTR(_CAST, 32643)
#define IDC_SIZEWE PTR(_CAST, 32644)
#define IDC_SIZENS PTR(_CAST, 32645)
#define IDC_SIZEALL PTR(_CAST, 32646)
#define IDC_NO PTR(_CAST, 32648)
#define IDC_APPSTARTING PTR(_CAST, 32650)
#define IDC_HELP PTR(_CAST, 32651)
#define IMAGE_BITMAP 0
#define IMAGE_ICON 1
#define IMAGE_CURSOR 2
#define IMAGE_ENHMETAFILE 3
#define BUTTON_IMAGELIST_ALIGN_BOTTOM 3
#define BUTTON_IMAGELIST_ALIGN_CENTER 4
#define BUTTON_IMAGELIST_ALIGN_LEFT 0
#define BUTTON_IMAGELIST_ALIGN_RIGHT 1
#define BUTTON_IMAGELIST_ALIGN_TOP 2
#define BCM_GETIDEALSIZE (BCM_FIRST + 0x0001)
#define BCM_GETIMAGELIST (BCM_FIRST + 0x0003)
#define BCM_SETIMAGELIST (BCM_FIRST + 0x0002)
#define LR_DEFAULTCOLOR 0x0000
#define LR_MONOCHROME 0x0001
#define LR_COLOR 0x0002
#define LR_COPYRETURNORG 0x0004
#define LR_COPYDELETEORG 0x0008
#define LR_LOADFROMFILE 0x0010
#define LR_LOADTRANSPARENT 0x0020
#define LR_DEFAULTSIZE 0x0040
#define LR_LOADREALSIZE 0x0080
#define LR_LOADMAP3DCOLORS 0x1000
#define LR_CREATEDIBSECTION 0x2000
#define LR_COPYFROMRESOURCE 0x4000
#define LR_SHARED 0x8000
#define DI_MASK 0x0001
#define DI_IMAGE 0x0002
#define DI_NORMAL 0x0003
#define DI_COMPAT 0x0004
#define DI_DEFAULTSIZE 0x0008
#define DI_NOMIRROR 0x0010
#define RES_ICON 1
#define RES_CURSOR 2
#define OBM_CLOSE 32754
#define OBM_UPARROW 32753
#define OBM_DNARROW 32752
#define OBM_RGARROW 32751
#define OBM_LFARROW 32750
#define OBM_REDUCE 32749
#define OBM_ZOOM 32748
#define OBM_RESTORE 32747
#define OBM_REDUCED 32746
#define OBM_ZOOMD 32745
#define OBM_RESTORED 32744
#define OBM_UPARROWD 32743
#define OBM_DNARROWD 32742
#define OBM_RGARROWD 32741
#define OBM_LFARROWD 32740
#define OBM_MNARROW 32739
#define OBM_COMBO 32738
#define OBM_UPARROWI 32737
#define OBM_DNARROWI 32736
#define OBM_RGARROWI 32735
#define OBM_LFARROWI 32734
#define OBM_OLD_CLOSE 32767
#define OBM_SIZE 32766
#define OBM_OLD_UPARROW 32765
#define OBM_OLD_DNARROW 32764
#define OBM_OLD_RGARROW 32763
#define OBM_OLD_LFARROW 32762
#define OBM_BTSIZE 32761
#define OBM_CHECK 32760
#define OBM_CHECKBOXES 32759
#define OBM_BTNCORNERS 32758
#define OBM_OLD_REDUCE 32757
#define OBM_OLD_ZOOM 32756
#define OBM_OLD_RESTORE 32755
#define OCR_NORMAL 32512
#define OCR_IBEAM 32513
#define OCR_WAIT 32514
#define OCR_CROSS 32515
#define OCR_UP 32516
#define OCR_SIZE 32640
#define OCR_ICON 32641
#define OCR_SIZENWSE 32642
#define OCR_SIZENESW 32643
#define OCR_SIZEWE 32644
#define OCR_SIZENS 32645
#define OCR_SIZEALL 32646
#define OCR_ICOCUR 32647
#define OCR_NO 32648
#define OCR_APPSTARTING 32650
#define OCR_HAND 32649
#define IDC_HAND PTR(_CAST, 32649)
#define OIC_SAMPLE 32512
#define OIC_HAND 32513
#define OIC_QUES 32514
#define OIC_BANG 32515
#define OIC_NOTE 32516
#define OIC_WINLOGO 32517
#define OIC_WARNING OIC_BANG
#define OIC_ERROR OIC_HAND
#define OIC_INFORMATION OIC_NOTE
#define ORD_LANGDRIVER 1
#define IDI_APPLICATION PTR(_CAST, 32512)
#define IDI_HAND PTR(_CAST, 32513)
#define IDI_QUESTION PTR(_CAST, 32514)
#define IDI_EXCLAMATION PTR(_CAST, 32515)
#define IDI_ASTERISK PTR(_CAST, 32516)
#define IDI_WINLOGO PTR(_CAST, 32517)
#define IDI_WARNING IDI_EXCLAMATION
#define IDI_ERROR IDI_HAND
#define IDI_INFORMATION IDI_ASTERISK
#define IDOK 1
#define IDCANCEL 2
#define IDABORT 3
#define IDRETRY 4
#define IDIGNORE 5
#define IDYES 6
#define IDNO 7
#define IDCLOSE 8
#define IDHELP 9
#define IDTRYAGAIN 10
#define IDCONTINUE 11
#define IDTIMEOUT 32000
#define ES_LEFT 0x0000L
#define ES_CENTER 0x0001L
#define ES_RIGHT 0x0002L
#define ES_MULTILINE 0x0004L
#define ES_UPPERCASE 0x0008L
#define ES_LOWERCASE 0x0010L
#define ES_PASSWORD 0x0020L
#define ES_AUTOVSCROLL 0x0040L
#define ES_AUTOHSCROLL 0x0080L
#define ES_NOHIDESEL 0x0100L
#define ES_OEMCONVERT 0x0400L
#define ES_READONLY 0x0800L
#define ES_WANTRETURN 0x1000L
#define ES_NUMBER 0x2000L
#define EN_SETFOCUS 0x0100
#define EN_KILLFOCUS 0x0200
#define EN_CHANGE 0x0300
#define EN_UPDATE 0x0400
#define EN_ERRSPACE 0x0500
#define EN_MAXTEXT 0x0501
#define EN_HSCROLL 0x0601
#define EN_VSCROLL 0x0602
#define EN_ALIGN_LTR_EC 0x0700
#define EN_ALIGN_RTL_EC 0x0701
#define EC_LEFTMARGIN 0x0001
#define EC_RIGHTMARGIN 0x0002
#define EC_USEFONTINFO 0xffff
#define EMSIS_COMPOSITIONSTRING 0x0001
#define EIMES_GETCOMPSTRATONCE 0x0001
#define EIMES_CANCELCOMPSTRINFOCUS 0x0002
#define EIMES_COMPLETECOMPSTRKILLFOCUS 0x0004
#define EM_GETSEL 0x00B0
#define EM_SETSEL 0x00B1
#define EM_GETRECT 0x00B2
#define EM_SETRECT 0x00B3
#define EM_SETRECTNP 0x00B4
#define EM_SCROLL 0x00B5
#define EM_LINESCROLL 0x00B6
#define EM_SCROLLCARET 0x00B7
#define EM_GETMODIFY 0x00B8
#define EM_SETMODIFY 0x00B9
#define EM_GETLINECOUNT 0x00BA
#define EM_LINEINDEX 0x00BB
#define EM_SETHANDLE 0x00BC
#define EM_GETHANDLE 0x00BD
#define EM_GETTHUMB 0x00BE
#define EM_LINELENGTH 0x00C1
#define EM_REPLACESEL 0x00C2
#define EM_GETLINE 0x00C4
#define EM_LIMITTEXT 0x00C5
#define EM_CANUNDO 0x00C6
#define EM_UNDO 0x00C7
#define EM_FMTLINES 0x00C8
#define EM_LINEFROMCHAR 0x00C9
#define EM_SETTABSTOPS 0x00CB
#define EM_SETPASSWORDCHAR 0x00CC
#define EM_EMPTYUNDOBUFFER 0x00CD
#define EM_GETFIRSTVISIBLELINE 0x00CE
#define EM_SETREADONLY 0x00CF
#define EM_SETWORDBREAKPROC 0x00D0
#define EM_GETWORDBREAKPROC 0x00D1
#define EM_GETPASSWORDCHAR 0x00D2
#define EM_SETMARGINS 0x00D3
#define EM_GETMARGINS 0x00D4
#define EM_SETLIMITTEXT EM_LIMITTEXT
#define EM_GETLIMITTEXT 0x00D5
#define EM_POSFROMCHAR 0x00D6
#define EM_CHARFROMPOS 0x00D7
#define EM_SETIMESTATUS 0x00D8
#define EM_GETIMESTATUS 0x00D9
#define WB_LEFT 0
#define WB_RIGHT 1
#define WB_ISDELIMITER 2
#define BS_PUSHBUTTON 0x00000000L
#define BS_DEFPUSHBUTTON 0x00000001L
#define BS_CHECKBOX 0x00000002L
#define BS_AUTOCHECKBOX 0x00000003L
#define BS_RADIOBUTTON 0x00000004L
#define BS_3STATE 0x00000005L
#define BS_AUTO3STATE 0x00000006L
#define BS_GROUPBOX 0x00000007L
#define BS_USERBUTTON 0x00000008L
#define BS_AUTORADIOBUTTON 0x00000009L
#define BS_PUSHBOX 0x0000000AL
#define BS_OWNERDRAW 0x0000000BL
#define BS_TYPEMASK 0x0000000FL
#define BS_LEFTTEXT 0x00000020L
#define BS_TEXT 0x00000000L
#define BS_ICON 0x00000040L
#define BS_BITMAP 0x00000080L
#define BS_LEFT 0x00000100L
#define BS_RIGHT 0x00000200L
#define BS_CENTER 0x00000300L
#define BS_TOP 0x00000400L
#define BS_BOTTOM 0x00000800L
#define BS_VCENTER 0x00000C00L
#define BS_PUSHLIKE 0x00001000L
#define BS_MULTILINE 0x00002000L
#define BS_NOTIFY 0x00004000L
#define BS_FLAT 0x00008000L
#define BS_RIGHTBUTTON BS_LEFTTEXT
#define BN_CLICKED 0
#define BN_PAINT 1
#define BN_HILITE 2
#define BN_UNHILITE 3
#define BN_DISABLE 4
#define BN_DOUBLECLICKED 5
#define BN_PUSHED BN_HILITE
#define BN_UNPUSHED BN_UNHILITE
#define BN_DBLCLK BN_DOUBLECLICKED
#define BN_SETFOCUS 6
#define BN_KILLFOCUS 7
#define BM_GETCHECK 0x00F0
#define BM_SETCHECK 0x00F1
#define BM_GETSTATE 0x00F2
#define BM_SETSTATE 0x00F3
#define BM_SETSTYLE 0x00F4
#define BM_CLICK 0x00F5
#define BM_GETIMAGE 0x00F6
#define BM_SETIMAGE 0x00F7
#define BST_UNCHECKED 0x0000
#define BST_CHECKED 0x0001
#define BST_INDETERMINATE 0x0002
#define BST_PUSHED 0x0004
#define BST_FOCUS 0x0008
#define SS_LEFT 0x00000000L
#define SS_CENTER 0x00000001L
#define SS_RIGHT 0x00000002L
#define SS_ICON 0x00000003L
#define SS_BLACKRECT 0x00000004L
#define SS_GRAYRECT 0x00000005L
#define SS_WHITERECT 0x00000006L
#define SS_BLACKFRAME 0x00000007L
#define SS_GRAYFRAME 0x00000008L
#define SS_WHITEFRAME 0x00000009L
#define SS_USERITEM 0x0000000AL
#define SS_SIMPLE 0x0000000BL
#define SS_LEFTNOWORDWRAP 0x0000000CL
#define SS_OWNERDRAW 0x0000000DL
#define SS_BITMAP 0x0000000EL
#define SS_ENHMETAFILE 0x0000000FL
#define SS_ETCHEDHORZ 0x00000010L
#define SS_ETCHEDVERT 0x00000011L
#define SS_ETCHEDFRAME 0x00000012L
#define SS_TYPEMASK 0x0000001FL
#define SS_REALSIZECONTROL 0x00000040L
#define SS_NOPREFIX 0x00000080L
#define SS_NOTIFY 0x00000100L
#define SS_CENTERIMAGE 0x00000200L
#define SS_RIGHTJUST 0x00000400L
#define SS_REALSIZEIMAGE 0x00000800L
#define SS_SUNKEN 0x00001000L
#define SS_EDITCONTROL 0x00002000L
#define SS_ENDELLIPSIS 0x00004000L
#define SS_PATHELLIPSIS 0x00008000L
#define SS_WORDELLIPSIS 0x0000C000L
#define SS_ELLIPSISMASK 0x0000C000L
#define STM_SETICON 0x0170
#define STM_GETICON 0x0171
#define STM_SETIMAGE 0x0172
#define STM_GETIMAGE 0x0173
#define STN_CLICKED 0
#define STN_DBLCLK 1
#define STN_ENABLE 2
#define STN_DISABLE 3
#define STM_MSGMAX 0x0174
#define WC_DIALOG PTR(_CAST, 0X8002)
#define DWL_MSGRESULT 0
#define DWL_DLGPROC 4
#define DWL_USER 8
#define DDL_READWRITE 0x0000
#define DDL_READONLY 0x0001
#define DDL_HIDDEN 0x0002
#define DDL_SYSTEM 0x0004
#define DDL_DIRECTORY 0x0010
#define DDL_ARCHIVE 0x0020
#define DDL_POSTMSGS 0x2000
#define DDL_DRIVES 0x4000
#define DDL_EXCLUSIVE 0x8000
#define DS_ABSALIGN 0x01L
#define DS_SYSMODAL 0x02L
#define DS_LOCALEDIT 0x20L
#define DS_SETFONT 0x40L
#define DS_MODALFRAME 0x80L
#define DS_NOIDLEMSG 0x100L
#define DS_SETFOREGROUND 0x200L
#define DS_3DLOOK 0x0004L
#define DS_FIXEDSYS 0x0008L
#define DS_NOFAILCREATE 0x0010L
#define DS_CONTROL 0x0400L
#define DS_CENTER 0x0800L
#define DS_CENTERMOUSE 0x1000L
#define DS_CONTEXTHELP 0x2000L
#define DS_SHELLFONT DS_SETFONT | DS_FIXEDSYS
#define DS_USEPIXELS 0x8000L
#define DM_GETDEFID (WM_USER+0)
#define DM_SETDEFID (WM_USER+1)
#define DM_REPOSITION (WM_USER+2)
#define PSM_PAGEINFO (WM_USER+100)
#define PSM_SHEETINFO (WM_USER+101)
#define PSI_SETACTIVE 0x0001L
#define PSI_KILLACTIVE 0x0002L
#define PSI_APPLY 0x0003L
#define PSI_RESET 0x0004L
#define PSI_HASHELP 0x0005L
#define PSI_HELP 0x0006L
#define PSI_CHANGED 0x0001L
#define PSI_GUISTART 0x0002L
#define PSI_REBOOT 0x0003L
#define PSI_GETSIBLINGS 0x0004L
#define DC_HASDEFID 0x534B
#define DLGC_WANTARROWS 0x0001
#define DLGC_WANTTAB 0x0002
#define DLGC_WANTALLKEYS 0x0004
#define DLGC_WANTMESSAGE 0x0004
#define DLGC_HASSETSEL 0x0008
#define DLGC_DEFPUSHBUTTON 0x0010
#define DLGC_UNDEFPUSHBUTTON 0x0020
#define DLGC_RADIOBUTTON 0x0040
#define DLGC_WANTCHARS 0x0080
#define DLGC_STATIC 0x0100
#define DLGC_BUTTON 0x2000
#define LB_CTLCODE 0L
#define LB_OKAY 0
#define LB_ERR (-1)
#define LB_ERRSPACE (-2)
#define LBN_ERRSPACE (-2)
#define LBN_SELCHANGE 1
#define LBN_DBLCLK 2
#define LBN_SELCANCEL 3
#define LBN_SETFOCUS 4
#define LBN_KILLFOCUS 5
#define LB_ADDSTRING 0x0180
#define LB_INSERTSTRING 0x0181
#define LB_DELETESTRING 0x0182
#define LB_SELITEMRANGEEX 0x0183
#define LB_RESETCONTENT 0x0184
#define LB_SETSEL 0x0185
#define LB_SETCURSEL 0x0186
#define LB_GETSEL 0x0187
#define LB_GETCURSEL 0x0188
#define LB_GETTEXT 0x0189
#define LB_GETTEXTLEN 0x018A
#define LB_GETCOUNT 0x018B
#define LB_SELECTSTRING 0x018C
#define LB_DIR 0x018D
#define LB_GETTOPINDEX 0x018E
#define LB_FINDSTRING 0x018F
#define LB_GETSELCOUNT 0x0190
#define LB_GETSELITEMS 0x0191
#define LB_SETTABSTOPS 0x0192
#define LB_GETHORIZONTALEXTENT 0x0193
#define LB_SETHORIZONTALEXTENT 0x0194
#define LB_SETCOLUMNWIDTH 0x0195
#define LB_ADDFILE 0x0196
#define LB_SETTOPINDEX 0x0197
#define LB_GETITEMRECT 0x0198
#define LB_GETITEMDATA 0x0199
#define LB_SETITEMDATA 0x019A
#define LB_SELITEMRANGE 0x019B
#define LB_SETANCHORINDEX 0x019C
#define LB_GETANCHORINDEX 0x019D
#define LB_SETCARETINDEX 0x019E
#define LB_GETCARETINDEX 0x019F
#define LB_SETITEMHEIGHT 0x01A0
#define LB_GETITEMHEIGHT 0x01A1
#define LB_FINDSTRINGEXACT 0x01A2
#define LB_SETLOCALE 0x01A5
#define LB_GETLOCALE 0x01A6
#define LB_SETCOUNT 0x01A7
#define LB_INITSTORAGE 0x01A8
#define LB_ITEMFROMPOINT 0x01A9
#define LB_MULTIPLEADDSTRING 0x01B1
#define LB_GETLISTBOXINFO 0x01B2
#define LB_MSGMAX 0x01B2
#define LBS_NOTIFY 0x0001L
#define LBS_SORT 0x0002L
#define LBS_NOREDRAW 0x0004L
#define LBS_MULTIPLESEL 0x0008L
#define LBS_OWNERDRAWFIXED 0x0010L
#define LBS_OWNERDRAWVARIABLE 0x0020L
#define LBS_HASSTRINGS 0x0040L
#define LBS_USETABSTOPS 0x0080L
#define LBS_NOINTEGRALHEIGHT 0x0100L
#define LBS_MULTICOLUMN 0x0200L
#define LBS_WANTKEYBOARDINPUT 0x0400L
#define LBS_EXTENDEDSEL 0x0800L
#define LBS_DISABLENOSCROLL 0x1000L
#define LBS_NODATA 0x2000L
#define LBS_NOSEL 0x4000L
#define LBS_COMBOBOX 0x8000L
#define LBS_STANDARD (LBS_NOTIFY | LBS_SORT | WS_VSCROLL | WS_BORDER)
#define CB_OKAY 0
#define CB_ERR (-1)
#define CB_ERRSPACE (-2)
#define CBN_ERRSPACE (-1)
#define CBN_SELCHANGE 1
#define CBN_DBLCLK 2
#define CBN_SETFOCUS 3
#define CBN_KILLFOCUS 4
#define CBN_EDITCHANGE 5
#define CBN_EDITUPDATE 6
#define CBN_DROPDOWN 7
#define CBN_CLOSEUP 8
#define CBN_SELENDOK 9
#define CBN_SELENDCANCEL 10
#define CBS_SIMPLE 0x0001L
#define CBS_DROPDOWN 0x0002L
#define CBS_DROPDOWNLIST 0x0003L
#define CBS_OWNERDRAWFIXED 0x0010L
#define CBS_OWNERDRAWVARIABLE 0x0020L
#define CBS_AUTOHSCROLL 0x0040L
#define CBS_OEMCONVERT 0x0080L
#define CBS_SORT 0x0100L
#define CBS_HASSTRINGS 0x0200L
#define CBS_NOINTEGRALHEIGHT 0x0400L
#define CBS_DISABLENOSCROLL 0x0800L
#define CBS_UPPERCASE 0x2000L
#define CBS_LOWERCASE 0x4000L
#define CB_GETEDITSEL 0x0140
#define CB_LIMITTEXT 0x0141
#define CB_SETEDITSEL 0x0142
#define CB_ADDSTRING 0x0143
#define CB_DIR 0x0145
#define CB_GETCOUNT 0x0146
#define CB_GETCURSEL 0x0147
#define CB_GETLBTEXT 0x0148
#define CB_GETLBTEXTLEN 0x0149
#define CB_INSERTSTRING 0x014A
#define CB_RESETCONTENT 0x014B
#define CB_FINDSTRING 0x014C
#define CB_SELECTSTRING 0x014D
#define CB_SETCURSEL 0x014E
#define CB_SHOWDROPDOWN 0x014F
#define CB_GETITEMDATA 0x0150
#define CB_SETITEMDATA 0x0151
#define CB_GETDROPPEDCONTROLRECT 0x0152
#define CB_SETITEMHEIGHT 0x0153
#define CB_GETITEMHEIGHT 0x0154
#define CB_SETEXTENDEDUI 0x0155
#define CB_GETEXTENDEDUI 0x0156
#define CB_GETDROPPEDSTATE 0x0157
#define CB_FINDSTRINGEXACT 0x0158
#define CB_SETLOCALE 0x0159
#define CB_GETLOCALE 0x015A
#define CB_GETTOPINDEX 0x015b
#define CB_SETTOPINDEX 0x015c
#define CB_GETHORIZONTALEXTENT 0x015d
#define CB_SETHORIZONTALEXTENT 0x015e
#define CB_GETDROPPEDWIDTH 0x015f
#define CB_SETDROPPEDWIDTH 0x0160
#define CB_INITSTORAGE 0x0161
#define CB_MULTIPLEADDSTRING 0x0163U
#define CB_GETCOMBOBOXINFO 0x0164
#define CB_MSGMAX 0x0164
#define SBS_HORZ 0x0000L
#define SBS_VERT 0x0001L
#define SBS_TOPALIGN 0x0002L
#define SBS_LEFTALIGN 0x0002L
#define SBS_BOTTOMALIGN 0x0004L
#define SBS_RIGHTALIGN 0x0004L
#define SBS_SIZEBOXTOPLEFTALIGN 0x0002L
#define SBS_SIZEBOXBOTTOMRIGHTALIGN 0x0004L
#define SBS_SIZEBOX 0x0008L
#define SBS_SIZEGRIP 0x0010L
#define SBM_SETPOS 0x00E0
#define SBM_GETPOS 0x00E1
#define SBM_SETRANGE 0x00E2
#define SBM_SETRANGEREDRAW 0x00E6
#define SBM_GETRANGE 0x00E3
#define SBM_ENABLE_ARROWS 0x00E4
#define SBM_SETSCROLLINFO 0x00E9
#define SBM_GETSCROLLINFO 0x00EA
#define SBM_GETSCROLLBARINFO 0x00EB
#define SIF_RANGE 0x0001
#define SIF_PAGE 0x0002
#define SIF_POS 0x0004
#define SIF_DISABLENOSCROLL 0x0008
#define SIF_TRACKPOS 0x0010
#define SIF_ALL (SIF_RANGE | SIF_PAGE | SIF_POS | SIF_TRACKPOS)
#define MDIS_ALLCHILDSTYLES 0x0001
#define MDITILE_VERTICAL 0x0000
#define MDITILE_HORIZONTAL 0x0001
#define MDITILE_SKIPDISABLED 0x0002
#define MDITILE_ZORDER 0x0004
#define IMC_GETCANDIDATEPOS 0x0007
#define IMC_SETCANDIDATEPOS 0x0008
#define IMC_GETCOMPOSITIONFONT 0x0009
#define IMC_SETCOMPOSITIONFONT 0x000A
#define IMC_GETCOMPOSITIONWINDOW 0x000B
#define IMC_SETCOMPOSITIONWINDOW 0x000C
#define IMC_GETSTATUSWINDOWPOS 0x000F
#define IMC_SETSTATUSWINDOWPOS 0x0010
#define IMC_CLOSESTATUSWINDOW 0x0021
#define IMC_OPENSTATUSWINDOW 0x0022
#define IMN_CLOSESTATUSWINDOW 0x0001
#define IMN_OPENSTATUSWINDOW 0x0002
#define IMN_CHANGECANDIDATE 0x0003
#define IMN_CLOSECANDIDATE 0x0004
#define IMN_OPENCANDIDATE 0x0005
#define IMN_SETCONVERSIONMODE 0x0006
#define IMN_SETSENTENCEMODE 0x0007
#define IMN_SETOPENSTATUS 0x0008
#define IMN_SETCANDIDATEPOS 0x0009
#define IMN_SETCOMPOSITIONFONT 0x000A
#define IMN_SETCOMPOSITIONWINDOW 0x000B
#define IMN_SETSTATUSWINDOWPOS 0x000C
#define IMN_GUIDELINE 0x000D
#define IMN_PRIVATE 0x000E
#define HELP_CONTEXT 0x0001L
#define HELP_QUIT 0x0002L
#define HELP_INDEX 0x0003L
#define HELP_CONTENTS 0x0003L
#define HELP_HELPONHELP 0x0004L
#define HELP_SETINDEX 0x0005L
#define HELP_SETCONTENTS 0x0005L
#define HELP_CONTEXTPOPUP 0x0008L
#define HELP_FORCEFILE 0x0009L
#define HELP_KEY 0x0101L
#define HELP_COMMAND 0x0102L
#define HELP_PARTIALKEY 0x0105L
#define HELP_MULTIKEY 0x0201L
#define HELP_SETWINPOS 0x0203L
#define HELP_CONTEXTMENU 0x000a
#define HELP_FINDER 0x000b
#define HELP_WM_HELP 0x000c
#define HELP_SETPOPUP_POS 0x000d
#define HELP_TCARD 0x8000
#define HELP_TCARD_DATA 0x0010
#define HELP_TCARD_OTHER_CALLER 0x0011
#define IDH_NO_HELP 28440
#define IDH_MISSING_CONTEXT 28441
#define IDH_GENERIC_HELP_BUTTON 28442
#define IDH_OK 28443
#define IDH_CANCEL 28444
#define IDH_HELP 28445
#define SPI_GETBEEP 1
#define SPI_SETBEEP 2
#define SPI_GETMOUSE 3
#define SPI_SETMOUSE 4
#define SPI_GETBORDER 5
#define SPI_SETBORDER 6
#define SPI_GETKEYBOARDSPEED 10
#define SPI_SETKEYBOARDSPEED 11
#define SPI_LANGDRIVER 12
#define SPI_ICONHORIZONTALSPACING 13
#define SPI_GETSCREENSAVETIMEOUT 14
#define SPI_SETSCREENSAVETIMEOUT 15
#define SPI_GETSCREENSAVEACTIVE 16
#define SPI_SETSCREENSAVEACTIVE 17
#define SPI_GETGRIDGRANULARITY 18
#define SPI_SETGRIDGRANULARITY 19
#define SPI_SETDESKWALLPAPER 20
#define SPI_SETDESKPATTERN 21
#define SPI_GETKEYBOARDDELAY 22
#define SPI_SETKEYBOARDDELAY 23
#define SPI_ICONVERTICALSPACING 24
#define SPI_GETICONTITLEWRAP 25
#define SPI_SETICONTITLEWRAP 26
#define SPI_GETMENUDROPALIGNMENT 27
#define SPI_SETMENUDROPALIGNMENT 28
#define SPI_SETDOUBLECLKWIDTH 29
#define SPI_SETDOUBLECLKHEIGHT 30
#define SPI_GETICONTITLELOGFONT 31
#define SPI_SETDOUBLECLICKTIME 32
#define SPI_SETMOUSEBUTTONSWAP 33
#define SPI_SETICONTITLELOGFONT 34
#define SPI_GETFASTTASKSWITCH 35
#define SPI_SETFASTTASKSWITCH 36
#define SPI_SETDRAGFULLWINDOWS 37
#define SPI_GETDRAGFULLWINDOWS 38
#define SPI_GETNONCLIENTMETRICS 41
#define SPI_SETNONCLIENTMETRICS 42
#define SPI_GETMINIMIZEDMETRICS 43
#define SPI_SETMINIMIZEDMETRICS 44
#define SPI_GETICONMETRICS 45
#define SPI_SETICONMETRICS 46
#define SPI_SETWORKAREA 47
#define SPI_GETWORKAREA 48
#define SPI_SETPENWINDOWS 49
#define SPI_GETHIGHCONTRAST 66
#define SPI_SETHIGHCONTRAST 67
#define SPI_GETKEYBOARDPREF 68
#define SPI_SETKEYBOARDPREF 69
#define SPI_GETSCREENREADER 70
#define SPI_SETSCREENREADER 71
#define SPI_GETANIMATION 72
#define SPI_SETANIMATION 73
#define SPI_GETFONTSMOOTHING 74
#define SPI_SETFONTSMOOTHING 75
#define SPI_SETDRAGWIDTH 76
#define SPI_SETDRAGHEIGHT 77
#define SPI_SETHANDHELD 78
#define SPI_GETLOWPOWERTIMEOUT 79
#define SPI_GETPOWEROFFTIMEOUT 80
#define SPI_SETLOWPOWERTIMEOUT 81
#define SPI_SETPOWEROFFTIMEOUT 82
#define SPI_GETLOWPOWERACTIVE 83
#define SPI_GETPOWEROFFACTIVE 84
#define SPI_SETLOWPOWERACTIVE 85
#define SPI_SETPOWEROFFACTIVE 86
#define SPI_SETCURSORS 87
#define SPI_SETICONS 88
#define SPI_GETDEFAULTINPUTLANG 89
#define SPI_SETDEFAULTINPUTLANG 90
#define SPI_SETLANGTOGGLE 91
#define SPI_GETWINDOWSEXTENSION 92
#define SPI_SETMOUSETRAILS 93
#define SPI_GETMOUSETRAILS 94
#define SPI_SETSCREENSAVERRUNNING 0x0061
#define SPI_SCREENSAVERRUNNING SPI_SETSCREENSAVERRUNNING
#define SPI_GETFILTERKEYS 50
#define SPI_SETFILTERKEYS 51
#define SPI_GETTOGGLEKEYS 52
#define SPI_SETTOGGLEKEYS 53
#define SPI_GETMOUSEKEYS 54
#define SPI_SETMOUSEKEYS 55
#define SPI_GETSHOWSOUNDS 56
#define SPI_SETSHOWSOUNDS 57
#define SPI_GETSTICKYKEYS 58
#define SPI_SETSTICKYKEYS 59
#define SPI_GETACCESSTIMEOUT 60
#define SPI_SETACCESSTIMEOUT 61
#define SPI_GETSERIALKEYS 62
#define SPI_SETSERIALKEYS 63
#define SPI_GETSOUNDSENTRY 64
#define SPI_SETSOUNDSENTRY 65
#define SPI_GETSNAPTODEFBUTTON 0x005F
#define SPI_SETSNAPTODEFBUTTON 0x0060
#define SPI_GETMOUSEHOVERWIDTH 0x0062
#define SPI_SETMOUSEHOVERWIDTH 0x0063
#define SPI_GETMOUSEHOVERHEIGHT 0x0064
#define SPI_SETMOUSEHOVERHEIGHT 0x0065
#define SPI_GETMOUSEHOVERTIME 0x0066
#define SPI_SETMOUSEHOVERTIME 0x0067
#define SPI_GETWHEELSCROLLLINES 0x0068
#define SPI_SETWHEELSCROLLLINES 0x0069
#define SPI_GETMENUSHOWDELAY 0x006A
#define SPI_SETMENUSHOWDELAY 0x006B
#define SPI_GETSHOWIMEUI 0x006E
#define SPI_SETSHOWIMEUI 0x006F
#define SPI_GETMOUSESPEED 0x0070
#define SPI_SETMOUSESPEED 0x0071
#define SPI_GETSCREENSAVERRUNNING 0x0072
#define SPI_GETDESKWALLPAPER 0x0073
#define SPI_GETACTIVEWINDOWTRACKING 0x1000
#define SPI_SETACTIVEWINDOWTRACKING 0x1001
#define SPI_GETMENUANIMATION 0x1002
#define SPI_SETMENUANIMATION 0x1003
#define SPI_GETCOMBOBOXANIMATION 0x1004
#define SPI_SETCOMBOBOXANIMATION 0x1005
#define SPI_GETLISTBOXSMOOTHSCROLLING 0x1006
#define SPI_SETLISTBOXSMOOTHSCROLLING 0x1007
#define SPI_GETGRADIENTCAPTIONS 0x1008
#define SPI_SETGRADIENTCAPTIONS 0x1009
#define SPI_GETKEYBOARDCUES 0x100A
#define SPI_SETKEYBOARDCUES 0x100B
#define SPI_GETMENUUNDERLINES SPI_GETKEYBOARDCUES
#define SPI_SETMENUUNDERLINES SPI_SETKEYBOARDCUES
#define SPI_GETACTIVEWNDTRKZORDER 0x100C
#define SPI_SETACTIVEWNDTRKZORDER 0x100D
#define SPI_GETHOTTRACKING 0x100E
#define SPI_SETHOTTRACKING 0x100F
#define SPI_GETMENUFADE 0x1012
#define SPI_SETMENUFADE 0x1013
#define SPI_GETSELECTIONFADE 0x1014
#define SPI_SETSELECTIONFADE 0x1015
#define SPI_GETTOOLTIPANIMATION 0x1016
#define SPI_SETTOOLTIPANIMATION 0x1017
#define SPI_GETTOOLTIPFADE 0x1018
#define SPI_SETTOOLTIPFADE 0x1019
#define SPI_GETCURSORSHADOW 0x101A
#define SPI_SETCURSORSHADOW 0x101B
#define SPI_GETMOUSESONAR 0x101C
#define SPI_SETMOUSESONAR 0x101D
#define SPI_GETMOUSECLICKLOCK 0x101E
#define SPI_SETMOUSECLICKLOCK 0x101F
#define SPI_GETMOUSEVANISH 0x1020
#define SPI_SETMOUSEVANISH 0x1021
#define SPI_GETFLATMENU 0x1022
#define SPI_SETFLATMENU 0x1023
#define SPI_GETDROPSHADOW 0x1024
#define SPI_SETDROPSHADOW 0x1025
#define SPI_GETBLOCKSENDINPUTRESETS 0x1026
#define SPI_SETBLOCKSENDINPUTRESETS 0x1027
#define SPI_GETUIEFFECTS 0x103E
#define SPI_SETUIEFFECTS 0x103F
#define SPI_GETFOREGROUNDLOCKTIMEOUT 0x2000
#define SPI_SETFOREGROUNDLOCKTIMEOUT 0x2001
#define SPI_GETACTIVEWNDTRKTIMEOUT 0x2002
#define SPI_SETACTIVEWNDTRKTIMEOUT 0x2003
#define SPI_GETFOREGROUNDFLASHCOUNT 0x2004
#define SPI_SETFOREGROUNDFLASHCOUNT 0x2005
#define SPI_GETCARETWIDTH 0x2006
#define SPI_SETCARETWIDTH 0x2007
#define SPI_GETMOUSECLICKLOCKTIME 0x2008
#define SPI_SETMOUSECLICKLOCKTIME 0x2009
#define SPI_GETFONTSMOOTHINGTYPE 0x200A
#define SPI_SETFONTSMOOTHINGTYPE 0x200B
#define FE_FONTSMOOTHINGSTANDARD 0x0001
#define FE_FONTSMOOTHINGCLEARTYPE 0x0002
#define FE_FONTSMOOTHINGDOCKING 0x8000
#define SPI_GETFONTSMOOTHINGCONTRAST 0x200C
#define SPI_SETFONTSMOOTHINGCONTRAST 0x200D
#define SPI_GETFOCUSBORDERWIDTH 0x200E
#define SPI_SETFOCUSBORDERWIDTH 0x200F
#define SPI_GETFOCUSBORDERHEIGHT 0x2010
#define SPI_SETFOCUSBORDERHEIGHT 0x2011
#define SPI_GETFONTSMOOTHINGORIENTATION 0x2012
#define SPI_SETFONTSMOOTHINGORIENTATION 0x2013
#define FE_FONTSMOOTHINGORIENTATIONBGR 0x0000
#define FE_FONTSMOOTHINGORIENTATIONRGB 0x0001
#define SPIF_UPDATEINIFILE 0x0001
#define SPIF_SENDWININICHANGE 0x0002
#define SPIF_SENDCHANGE SPIF_SENDWININICHANGE
#define METRICS_USEDEFAULT -1
#define ARW_BOTTOMLEFT 0x0000L
#define ARW_BOTTOMRIGHT 0x0001L
#define ARW_TOPLEFT 0x0002L
#define ARW_TOPRIGHT 0x0003L
#define ARW_STARTMASK 0x0003L
#define ARW_STARTRIGHT 0x0001L
#define ARW_STARTTOP 0x0002L
#define ARW_LEFT 0x0000L
#define ARW_RIGHT 0x0000L
#define ARW_UP 0x0004L
#define ARW_DOWN 0x0004L
#define ARW_HIDE 0x0008L
#define ARW_VALID 0x000FL
#define SERKF_SERIALKEYSON 0x00000001
#define SERKF_AVAILABLE 0x00000002
#define SERKF_INDICATOR 0x00000004
#define HCF_HIGHCONTRASTON 0x00000001
#define HCF_AVAILABLE 0x00000002
#define HCF_HOTKEYACTIVE 0x00000004
#define HCF_CONFIRMHOTKEY 0x00000008
#define HCF_HOTKEYSOUND 0x00000010
#define HCF_INDICATOR 0x00000020
#define HCF_HOTKEYAVAILABLE 0x00000040
#define HCF_LOGONDESKTOP 0x00000100
#define HCF_DEFAULTDESKTOP 0x00000200
#define CDS_UPDATEREGISTRY 0x00000001
#define CDS_TEST 0x00000002
#define CDS_FULLSCREEN 0x00000004
#define CDS_GLOBAL 0x00000008
#define CDS_SET_PRIMARY 0x00000010
#define CDS_VIDEOPARAMETERS 0x00000020
#define CDS_RESET 0x40000000
#define CDS_NORESET 0x10000000
#define DISP_CHANGE_SUCCESSFUL 0
#define DISP_CHANGE_RESTART 1
#define DISP_CHANGE_FAILED -1
#define DISP_CHANGE_BADMODE -2
#define DISP_CHANGE_NOTUPDATED -3
#define DISP_CHANGE_BADFLAGS -4
#define DISP_CHANGE_BADPARAM -5
#define DISP_CHANGE_BADDUALVIEW -6
#define ENUM_CURRENT_SETTINGS 0xFFFFFFFU
#define ENUM_REGISTRY_SETTINGS 0xFFFFFFEU
#define FKF_FILTERKEYSON 0x00000001
#define FKF_AVAILABLE 0x00000002
#define FKF_HOTKEYACTIVE 0x00000004
#define FKF_CONFIRMHOTKEY 0x00000008
#define FKF_HOTKEYSOUND 0x00000010
#define FKF_INDICATOR 0x00000020
#define FKF_CLICKON 0x00000040
#define SKF_STICKYKEYSON 0x00000001
#define SKF_AVAILABLE 0x00000002
#define SKF_HOTKEYACTIVE 0x00000004
#define SKF_CONFIRMHOTKEY 0x00000008
#define SKF_HOTKEYSOUND 0x00000010
#define SKF_INDICATOR 0x00000020
#define SKF_AUDIBLEFEEDBACK 0x00000040
#define SKF_TRISTATE 0x00000080
#define SKF_TWOKEYSOFF 0x00000100
#define SKF_LALTLATCHED 0x10000000
#define SKF_LCTLLATCHED 0x04000000
#define SKF_LSHIFTLATCHED 0x01000000
#define SKF_RALTLATCHED 0x20000000
#define SKF_RCTLLATCHED 0x08000000
#define SKF_RSHIFTLATCHED 0x02000000
#define SKF_LWINLATCHED 0x40000000
#define SKF_RWINLATCHED 0x80000000
#define SKF_LALTLOCKED 0x00100000
#define SKF_LCTLLOCKED 0x00040000
#define SKF_LSHIFTLOCKED 0x00010000
#define SKF_RALTLOCKED 0x00200000
#define SKF_RCTLLOCKED 0x00080000
#define SKF_RSHIFTLOCKED 0x00020000
#define SKF_LWINLOCKED 0x00400000
#define SKF_RWINLOCKED 0x00800000
#define MKF_MOUSEKEYSON 0x00000001
#define MKF_AVAILABLE 0x00000002
#define MKF_HOTKEYACTIVE 0x00000004
#define MKF_CONFIRMHOTKEY 0x00000008
#define MKF_HOTKEYSOUND 0x00000010
#define MKF_INDICATOR 0x00000020
#define MKF_MODIFIERS 0x00000040
#define MKF_REPLACENUMBERS 0x00000080
#define MKF_LEFTBUTTONSEL 0x10000000
#define MKF_RIGHTBUTTONSEL 0x20000000
#define MKF_LEFTBUTTONDOWN 0x01000000
#define MKF_RIGHTBUTTONDOWN 0x02000000
#define MKF_MOUSEMODE 0x80000000
#define ATF_TIMEOUTON 0x00000001
#define ATF_ONOFFFEEDBACK 0x00000002
#define SSGF_NONE 0
#define SSGF_DISPLAY 3
#define SSTF_NONE 0
#define SSTF_CHARS 1
#define SSTF_BORDER 2
#define SSTF_DISPLAY 3
#define SSWF_NONE 0
#define SSWF_TITLE 1
#define SSWF_WINDOW 2
#define SSWF_DISPLAY 3
#define SSWF_CUSTOM 4
#define SSF_SOUNDSENTRYON 0x00000001
#define SSF_AVAILABLE 0x00000002
#define SSF_INDICATOR 0x00000004
#define TKF_TOGGLEKEYSON 0x00000001
#define TKF_AVAILABLE 0x00000002
#define TKF_HOTKEYACTIVE 0x00000004
#define TKF_CONFIRMHOTKEY 0x00000008
#define TKF_HOTKEYSOUND 0x00000010
#define TKF_INDICATOR 0x00000020
#define SLE_ERROR 0x00000001
#define SLE_MINORERROR 0x00000002
#define SLE_WARNING 0x00000003
#define MONITOR_DEFAULTTONULL 0x00000000
#define MONITOR_DEFAULTTOPRIMARY 0x00000001
#define MONITOR_DEFAULTTONEAREST 0x00000002
#define CCHILDREN_TITLEBAR 5
#define CCHILDREN_SCROLLBAR 5
#define CCHILDREN_FRAME 7
#define OBJID_WINDOW 0x00000000L
#define OBJID_SYSMENU 0xFFFFFFFFL
#define OBJID_TITLEBAR 0xFFFFFFFEL
#define OBJID_MENU 0xFFFFFFFDL
#define OBJID_CLIENT 0xFFFFFFFCL
#define OBJID_VSCROLL 0xFFFFFFFBL
#define OBJID_HSCROLL 0xFFFFFFFAL
#define OBJID_SIZEGRIP 0xFFFFFFF9L
#define OBJID_CARET 0xFFFFFFF8L
#define OBJID_CURSOR 0xFFFFFFF7L
#define OBJID_ALERT 0xFFFFFFF6L
#define OBJID_SOUND 0xFFFFFFF5L
#define OBJID_QUERYCLASSNAMEIDX 0xFFFFFFF4L
#define OBJID_NATIVEOM 0xFFFFFFF0L
#define ASC_NUL 0x00
#define ASC_SOH 0x01
#define ASC_STX 0x02
#define ASC_ETX 0x03
#define ASC_EOT 0x04
#define ASC_ENQ 0x05
#define ASC_ACK 0x06
#define ASC_BEL 0x07
#define ASC_BS 0x08
#define ASC_HT 0x09
#define ASC_LF 0x0A
#define ASC_VT 0x0B
#define ASC_FF 0x0C
#define ASC_CR 0x0D
#define ASC_SO 0x0E
#define ASC_SI 0x0F
#define ASC_DLE 0x10
#define ASC_DC1 0x11
#define ASC_DC2 0x12
#define ASC_DC3 0x13
#define ASC_DC4 0x14
#define ASC_NAK 0x15
#define ASC_SYN 0x16
#define ASC_ETB 0x17
#define ASC_CAN 0x18
#define ASC_EM 0x19
#define ASC_SS 0x1A
#define ASC_ESC 0x1B
#define ASC_FS 0x1C
#define ASC_GS 0x1D
#define ASC_RS 0x1E
#define ASC_US 0x1F
#define ASC_SP 0x20
#define ASC_Exclamation 0x21
#define ASC_Quotation 0x22
#define ASC_DoubleQMark 0x22
#define ASC_Number 0x23
#define ASC_Dollar 0x24
#define ASC_Percent 0x25
#define ASC_Ampersand 0x26
#define ASC_Apostrophe 0x27
#define ASC_SingleQMark 0x27
#define ASC_LeftP 0x28
#define ASC_RightP 0x29
#define ASC_Asterisk 0x2A
#define ASC_Plus 0x2B
#define ASC_Comma 0x2C
#define ASC_Minus 0x2D
#define ASC_Hyphen 0x2D
#define ASC_Dot 0x2E
#define ASC_Period 0x2E
#define ASC_FullStop 0x2E
#define ASC_Solidus 0x2F
#define ASC_Slash 0x2F
#define ASC_0 0x30
#define ASC_1 0x31
#define ASC_2 0x32
#define ASC_3 0x33
#define ASC_4 0x34
#define ASC_5 0x35
#define ASC_6 0x36
#define ASC_7 0x37
#define ASC_8 0x38
#define ASC_9 0x39
#define ASC_Colon 0x3A
#define ASC_Semicolon 0x3B
#define ASC_Less 0x3C
#define ASC_Equals 0x3D
#define ASC_Greater 0x3E
#define ASC_Question 0x3F
#define ASC_AT 0x40
#define ASC_A 0x41
#define ASC_B 0x42
#define ASC_C 0x43
#define ASC_D 0x44
#define ASC_E 0x45
#define ASC_F 0x46
#define ASC_G 0x47
#define ASC_H 0x48
#define ASC_I 0x49
#define ASC_J 0x4A
#define ASC_K 0x4B
#define ASC_L 0x4C
#define ASC_M 0x4D
#define ASC_N 0x4E
#define ASC_O 0x4F
#define ASC_P 0x50
#define ASC_Q 0x51
#define ASC_R 0x52
#define ASC_S 0x53
#define ASC_T 0x54
#define ASC_U 0x55
#define ASC_V 0x56
#define ASC_W 0x57
#define ASC_X 0x58
#define ASC_Y 0x59
#define ASC_Z 0x5A
#define ASC_LeftSq 0x5B
#define ASC_BackSlash 0x5C
#define ASC_RightSq 0x5D
#define ASC_Circumflex 0x5E
#define ASC_Underscore 0x5f
#define ASC_a_ 0x61
#define ASC_b_ 0x62
#define ASC_c_ 0x63
#define ASC_d_ 0x64
#define ASC_e_ 0x65
#define ASC_f_ 0x66
#define ASC_g_ 0x67
#define ASC_h_ 0x68
#define ASC_i_ 0x69
#define ASC_j_ 0x6A
#define ASC_k_ 0x6B
#define ASC_l_ 0x6C
#define ASC_m_ 0x6D
#define ASC_n_ 0x6E
#define ASC_o_ 0x6F
#define ASC_p_ 0x70
#define ASC_q_ 0x71
#define ASC_r_ 0x72
#define ASC_s_ 0x73
#define ASC_t_ 0x74
#define ASC_u_ 0x75
#define ASC_v_ 0x76
#define ASC_w_ 0x77
#define ASC_x_ 0x78
#define ASC_y_ 0x79
#define ASC_z_ 0x7A
#define ASC_LeftCurly 0x7B
#define ASC_VertLine 0x7C
#define ASC_RightCurly 0x7D
#define ASC_Tilde 0x7E
#define ASC_Delete 0x7f
#define SIZEOFWIN95MENUITEMINFO 44
#define MIIM_STRING 0x00000040
#define MIIM_BITMAP 0x00000080
#define MIIM_FTYPE 0x00000100
#define EM_SETUNDOLIMIT (WM_USER + 82) 
#define EM_REDO (WM_USER + 84)
#define EM_CANREDO (WM_USER + 85)
#define EM_GETUNDONAME (WM_USER + 86)
#define EM_GETREDONAME (WM_USER + 87)
#define EM_STOPGROUPTYPING (WM_USER + 88)
#define EM_SETTEXTMODE (WM_USER + 89)
#define EM_GETTEXTMODE (WM_USER + 90)
#define TM_PLAINTEXT 1
#define TM_RICHTEXT 2 
#define TM_SINGLELEVELUNDO 4
#define TM_MULTILEVELUNDO 8 
#define TM_SINGLECODEPAGE 16
#define TM_MULTICODEPAGE 32 
#define EM_AUTOURLDETECT (WM_USER + 91)
#define EM_GETAUTOURLDETECT (WM_USER + 92)
#define EM_SETPALETTE (WM_USER + 93)
#define EM_GETTEXTEX (WM_USER + 94)
#define EM_GETTEXTLENGTHEX (WM_USER + 95)
#define STATE_SYSTEM_UNAVAILABLE 0x00000001U
#define STATE_SYSTEM_SELECTED 0x00000002U
#define STATE_SYSTEM_FOCUSED 0x00000004U
#define STATE_SYSTEM_PRESSED 0x00000008U
#define STATE_SYSTEM_CHECKED 0x00000010U
#define STATE_SYSTEM_MIXED 0x00000020U
#define STATE_SYSTEM_READONLY 0x00000040U
#define STATE_SYSTEM_HOTTRACKED 0x00000080U
#define STATE_SYSTEM_DEFAULT 0x00000100U
#define STATE_SYSTEM_EXPANDED 0x00000200U
#define STATE_SYSTEM_COLLAPSED 0x00000400U
#define STATE_SYSTEM_BUSY 0x00000800U
#define STATE_SYSTEM_FLOATING 0x00001000U
#define STATE_SYSTEM_MARQUEED 0x00002000U
#define STATE_SYSTEM_ANIMATED 0x00004000U
#define STATE_SYSTEM_INVISIBLE 0x00008000U
#define STATE_SYSTEM_OFFSCREEN 0x00010000U
#define STATE_SYSTEM_SIZEABLE 0x00020000U
#define STATE_SYSTEM_MOVEABLE 0x00040000U
#define STATE_SYSTEM_SELFVOICING 0x00080000U
#define STATE_SYSTEM_FOCUSABLE 0x00100000U
#define STATE_SYSTEM_SELECTABLE 0x00200000U
#define STATE_SYSTEM_LINKED 0x00400000U
#define STATE_SYSTEM_TRAVERSED 0x00800000U
#define STATE_SYSTEM_MULTISELECTABLE 0x01000000U
#define STATE_SYSTEM_EXTSELECTABLE 0x02000000U
#define STATE_SYSTEM_ALERT_LOW 0x04000000U
#define STATE_SYSTEM_ALERT_MEDIUM 0x08000000U
#define STATE_SYSTEM_ALERT_HIGH 0x10000000U
#define STATE_SYSTEM_VALID 0x1FFFFFFFU
#define VS_FILE_INFO RT_VERSION
#define VS_VERSION_INFO 1
#define VS_USER_DEFINED 100
#define VS_FFI_SIGNATURE 0xFEEF04BDL
#define VS_FFI_STRUCVERSION 0x00010000L
#define VS_FFI_FILEFLAGSMASK 0x0000003FL
#define VS_FF_DEBUG 0x00000001L
#define VS_FF_PRERELEASE 0x00000002L
#define VS_FF_PATCHED 0x00000004L
#define VS_FF_PRIVATEBUILD 0x00000008L
#define VS_FF_INFOINFERRED 0x00000010L
#define VS_FF_SPECIALBUILD 0x00000020L
#define VOS_UNKNOWN 0x00000000L
#define VOS_DOS 0x00010000L
#define VOS_OS216 0x00020000L
#define VOS_OS232 0x00030000L
#define VOS_NT 0x00040000L
#define VOS_WINCE 0x00050000L
#define VOS__BASE 0x00000000L
#define VOS__WINDOWS16 0x00000001L
#define VOS__PM16 0x00000002L
#define VOS__PM32 0x00000003L
#define VOS__WINDOWS32 0x00000004L
#define VOS_DOS_WINDOWS16 0x00010001L
#define VOS_DOS_WINDOWS32 0x00010004L
#define VOS_OS216_PM16 0x00020002L
#define VOS_OS232_PM32 0x00030003L
#define VOS_NT_WINDOWS32 0x00040004L
#define VFT_UNKNOWN 0x00000000L
#define VFT_APP 0x00000001L
#define VFT_DLL 0x00000002L
#define VFT_DRV 0x00000003L
#define VFT_FONT 0x00000004L
#define VFT_VXD 0x00000005L
#define VFT_STATIC_LIB 0x00000007L
#define VFT2_UNKNOWN 0x00000000L
#define VFT2_DRV_PRINTER 0x00000001L
#define VFT2_DRV_KEYBOARD 0x00000002L
#define VFT2_DRV_LANGUAGE 0x00000003L
#define VFT2_DRV_DISPLAY 0x00000004L
#define VFT2_DRV_MOUSE 0x00000005L
#define VFT2_DRV_NETWORK 0x00000006L
#define VFT2_DRV_SYSTEM 0x00000007L
#define VFT2_DRV_INSTALLABLE 0x00000008L
#define VFT2_DRV_SOUND 0x00000009L
#define VFT2_DRV_COMM 0x0000000AL
#define VFT2_DRV_INPUTMETHOD 0x0000000BL
#define VFT2_DRV_VERSIONED_PRINTER 0x0000000CL
#define VFT2_FONT_RASTER 0x00000001L
#define VFT2_FONT_VECTOR 0x00000002L
#define VFT2_FONT_TRUETYPE 0x00000003L
#define VFFF_ISSHAREDFILE 0x0001
#define VFF_CURNEDEST 0x0001
#define VFF_FILEINUSE 0x0002
#define VFF_BUFFTOOSMALL 0x0004
#define VIFF_FORCEINSTALL 0x0001
#define VIFF_DONTDELETEOLD 0x0002
#define VIF_TEMPFILE 0x00000001L
#define VIF_MISMATCH 0x00000002L
#define VIF_SRCOLD 0x00000004L
#define VIF_DIFFLANG 0x00000008L
#define VIF_DIFFCODEPG 0x00000010L
#define VIF_DIFFTYPE 0x00000020L
#define VIF_WRITEPROT 0x00000040L
#define VIF_FILEINUSE 0x00000080L
#define VIF_OUTOFSPACE 0x00000100L
#define VIF_ACCESSVIOLATION 0x00000200L
#define VIF_SHARINGVIOLATION 0x00000400L
#define VIF_CANNOTCREATE 0x00000800L
#define VIF_CANNOTDELETE 0x00001000L
#define VIF_CANNOTRENAME 0x00002000L
#define VIF_CANNOTDELETECUR 0x00004000L
#define VIF_OUTOFMEMORY 0x00008000L
#define VIF_CANNOTREADSRC 0x00010000L
#define VIF_CANNOTREADDST 0x00020000L
#define VIF_BUFFTOOSMALL 0x00040000L
#define VIF_CANNOTLOADLZ32 0x00080000L
#define VIF_CANNOTLOADCABINET 0x00100000L
#define MEMCTX_TASK 1
#define MEMCTX_SHARED 2
#define MEMCTX_MACSYSTEM 3
#define MEMCTX_UNKNOWN -1
#define MEMCTX_SAME -2
#define CLSCTX_INPROC_SERVER16 8
#define MSHLFLAGS_NORMAL 0
#define MSHLFLAGS_TABLESTRONG 1
#define MSHLFLAGS_TABLEWEAK 2
#define MSHCTX_LOCAL 0
#define MSHCTX_NOSHAREDMEM 1
#define MSHCTX_DIFFERENTMACHINE 2
#define MSHCTX_INPROC 3
#define DVASPECT_CONTENT 1
#define DVASPECT_THUMBNAIL 2
#define DVASPECT_ICON 4
#define DVASPECT_DOCPRINT 8
#define STGC_DEFAULT 0
#define STGC_OVERWRITE 1
#define STGC_ONLYIFCURRENT 2
#define STGC_DANGEROUSLYCOMMITMERELYTODISKCACHE 4
#define STGMOVE_MOVE 0
#define STGMOVE_COPY 1
#define STATFLAG_DEFAULT 0
#define STATFLAG_NONAME 1
