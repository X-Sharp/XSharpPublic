///////////////////////////////////////////////////////////////////////////
// VORDDClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// RDD Classes library
//

#define DBCCON TRUE
#define DBCCOFF FALSE
#define DBCCREADONLY FALSE
#define DBCCUPDATE TRUE
#define DBEXCLUSIVE FALSE
#define DBREADONLY TRUE
#define DBREADWRITE FALSE
#define DBSCOPEALL FALSE
#define DBSCOPEREST TRUE
#define DBSELECTIONEMPTY -2
#define DBSELECTIONBOF -1
#define DBSELECTIONEOF 1
#define DBSELECTIONFOUND 2
#define DBSELECTIONNULL 0
#define DBSHARED TRUE
#define ORD_KEYCOUNT 2
#define ORD_KEYDEC 4
#define ORD_KEYEXPR 3
#define ORD_KEYINFO 8
#define ORD_KEYSIZE 3
#define ORD_KEYTYPE 1
#define BUFFER_VALUE 1
#define BUFFER_BLOB_VALUE 2
#define BUFFER_IS_CHANGED 2
#define BUFFER_IS_BLOB 2
