///////////////////////////////////////////////////////////////////////////
// VOInternetServerClasses.vh
//
// Copyright (c) Grafx Database Systems, Inc.  All rights reserved.
//
// Vulcan.NET preprocessor directives for the Visual Objects-compatible
// Internet Server Classes library
//

#define MAX_BUFFER 256
#define CR _CHR(13)
#define LF _CHR(10)
#define HSE_IO_ASYNC 0x00000002
#define HSE_IO_DISCONNECT_AFTER_SEND 0x00000004
#define HSE_IO_SEND_HEADERS 0x00000008
#define HSE_IO_SYNC 0x00000001
#define HSE_LOG_BUFFER_LEN 80
#define HSE_MAX_EXT_DLL_NAME_LEN 256
#define HSE_REQ_BASE 0
#define HSE_REQ_DONE_WITH_SESSION ( HSE_REQ_BASE + 4 )
#define HSE_REQ_END_RESERVED 1000
#define HSE_REQ_GET_SSPI_INFO (HSE_REQ_END_RESERVED+2)
#define HSE_REQ_MAP_URL_TO_PATH (HSE_REQ_END_RESERVED+1)
#define HSE_REQ_SEND_RESPONSE_HEADER ( HSE_REQ_BASE + 3 )
#define HSE_REQ_SEND_URL ( HSE_REQ_BASE + 2 )
#define HSE_REQ_SEND_URL_EX (HSE_REQ_END_RESERVED+4)
#define HSE_REQ_SEND_URL_REDIRECT_RESP ( HSE_REQ_BASE + 1 )
#define HSE_APPEND_LOG_PARAMETER (HSE_REQ_END_RESERVED+3)
#define HSE_STATUS_ERROR 4
#define HSE_STATUS_PENDING 3
#define HSE_STATUS_SUCCESS 1
#define HSE_STATUS_SUCCESS_AND_KEEP_CONN 2
#define HSE_TERM_ADVISORY_UNLOAD 0x00000001
#define HSE_TERM_MUST_UNLOAD 0x00000002
#define HSE_VERSION_MAJOR 2
#define HSE_VERSION_MINOR 0
#define HTTP_FILTER_REVISION 2L
#define HTTP_GET "GET"
#define HTTP_POST "POST"
#define SF_DENIED_APPLICATION 0x00000008
#define SF_DENIED_BY_CONFIG 0x00010000
#define SF_DENIED_FILTER 0x00000004
#define SF_DENIED_LOGON 0x00000001
#define SF_DENIED_RESOURCE 0x00000002
#define SF_MAX_FILTER_DESC_LEN 257
#define SF_MAX_PASSWORD 257
#define SF_MAX_USERNAME 257
#define SF_NOTIFY_ACCESS_DENIED 0x00000800
#define SF_NOTIFY_AUTHENTICATION 0x00002000
#define SF_NOTIFY_END_OF_NET_SESSION 0x00000100
#define SF_NOTIFY_LOG 0x00000200
#define SF_NOTIFY_NONSECURE_PORT 0x00000002
#define SF_NOTIFY_ORDER_LOW 0x00020000
#define SF_NOTIFY_ORDER_DEFAULT SF_NOTIFY_ORDER_LOW
#define SF_NOTIFY_ORDER_HIGH 0x00080000
#define SF_NOTIFY_ORDER_MEDIUM 0x00040000
#define SF_NOTIFY_ORDER_MASK SF_NOTIFY_ORDER_HIGH + SF_NOTIFY_ORDER_MEDIUM + SF_NOTIFY_ORDER_LOW
#define SF_NOTIFY_PREPROC_HEADERS 0x00004000
#define SF_NOTIFY_READ_RAW_DATA 0x00008000
#define SF_NOTIFY_SECURE_PORT 0x00000001
#define SF_NOTIFY_SEND_RAW_DATA 0x00000400
#define SF_NOTIFY_URL_MAP 0x00001000
#define SF_REQ_ADD_HEADERS_ON_DENIAL 1
#define SF_REQ_SEND_RESPONSE_HEADER 0
#define SF_REQ_SET_NEXT_READ_SIZE 2
#define SF_REQ_SET_PROXY_INFO 3
#define SF_STATUS_REQ_ERROR 0x8000004
#define SF_STATUS_REQ_FINISHED 0x8000000
#define SF_STATUS_REQ_FINISHED_KEEP_CONN 0x8000001
#define SF_STATUS_REQ_HANDLED_NOTIFICATION 0x8000003
#define SF_STATUS_REQ_NEXT_NOTIFICATION 0x8000002
#define SF_STATUS_REQ_READ_NEXT 0x8000005
